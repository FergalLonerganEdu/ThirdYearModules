module lookuptable_rom_1 ( input [4:0]	addr,
						output [35:0]	data
					 );
				
	// ROM definition				
	parameter [0:27][35:0] ROM = {
   36'b000000000100000000000010000100000000, //p1
	36'b010000000000000000010000001000000000,
	36'b010010000100000000010010000100000010, //p2
	36'b000110000100000000000110000100001000,
	36'b000010010100000000000010010110000000,
	36'b000010000100010000100010000100010000,
	36'b000010000100000100001010000100000100,
	36'b000010000100000001100010000100000001,
	36'b000010000101000000000010100101000000,
	36'b010110000100000010010110000110000010, //p3
	36'b010010010100000010010010010110000010,
	36'b010010000100010010010010000110010010,
	36'b010010000100000110010010000110000110,
	36'b010010000101000010010010100101000010,
	36'b010110100101000010010110100101001010, //p4
	36'b010010100101000110001010100101000110,
	36'b010010100101010010011010100101010010,
	36'b010110000100001000010110000100001010, //p5
	36'b000110000100001001100110000100001001,
	36'b000110000100011000000110100100011000,
	36'b000110010100001000000110010110001000,
	36'b000110000101001000000110100101001000,
	36'b010110010100001010010110010110001010, //p6
	36'b010110000100011010010110000110011010,
	36'b010110000101001010010110000101101010,
	36'b100110010100001001100110010110001001, //p7
	36'b100110000101001001100110100101001001,
	36'b100110000100011001100110100100011001
};


assign data = ROM[addr];

endmodule  
