module shape_rom ( input [8:0]	addr,
						output [119:0]	data
					 );

	parameter ADDR_WIDTH = 9;
   parameter DATA_WIDTH =  120;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:359][DATA_WIDTH-1:0] ROM = {
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
         
// code x01
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
		  120'b000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000,
		  120'b000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000,
		  120'b000000000000000000000000000000000000000000011111111111111111111111111111111110000000000000000000000000000000000000000000,
		  120'b000000000000000000000000000000000000000011111111111111111111111111111111111111110000000000000000000000000000000000000000,
		  120'b000000000000000000000000000000000000001111111111111111111111111111111111111111111100000000000000000000000000000000000000,
		  120'b000000000000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000000000,
		  120'b000000000000000000000000000000000011111111111111111111111111111111111111111111111111110000000000000000000000000000000000,
		  120'b000000000000000000000000000000000111111111111111111111111111111111111111111111111111111000000000000000000000000000000000,
		  120'b000000000000000000000000000000011111111111111111111111111111111111111111111111111111111110000000000000000000000000000000,
		  120'b000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000,
		  120'b000000000000000000000000000001111111111111111111111000000000000000000111111111111111111111100000000000000000000000000000,
		  120'b000000000000000000000000000011111111111111111111000000000000000000000000111111111111111111110000000000000000000000000000,
		  120'b000000000000000000000000001111111111111111111000000000000000000000000000000111111111111111111100000000000000000000000000,
		  120'b000000000000000000000000011111111111111111100000000000000000000000000000000001111111111111111110000000000000000000000000,
		  120'b000000000000000000000000111111111111111110000000000000000000000000000000000000011111111111111111000000000000000000000000,
		  120'b000000000000000000000001111111111111111000000000000000000000000000000000000000000111111111111111100000000000000000000000,
		  120'b000000000000000000000011111111111111100000000000000000000000000000000000000000000001111111111111110000000000000000000000,
		  120'b000000000000000000000011111111111111000000000000000000000000000000000000000000000000111111111111110000000000000000000000,
		  120'b000000000000000000000111111111111110000000000000000000000000000000000000000000000000011111111111111000000000000000000000,
		  120'b000000000000000000001111111111111100000000000000000000000000000000000000000000000000001111111111111100000000000000000000,
		  120'b000000000000000000011111111111110000000000000000000000000000000000000000000000000000000011111111111110000000000000000000,
		  120'b000000000000000000011111111111100000000000000000000000000000000000000000000000000000000001111111111110000000000000000000,
		  120'b000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000,
		  120'b000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000,
		  120'b000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000,
		  120'b000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000,
		  120'b000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000000,
		  120'b000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000,
		  120'b000000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000,
		  120'b000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000000,
		  120'b000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000000,
		  120'b000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000,
		  120'b000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000,
		  120'b000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000,
		  120'b000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000,
		  120'b000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000,
		  120'b000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000,
		  120'b000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000,
		  120'b000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000,
		  120'b000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000,
		  120'b000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000,
		  120'b000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000,
		  120'b000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000,
		  120'b000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000,
		  120'b000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000,
		  120'b000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000,
		  120'b000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000,
		  120'b000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000,
		  120'b000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000,
		  120'b000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000,
		  120'b000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000,
		  120'b000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000,
		  120'b000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000,
		  120'b000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000,
		  120'b000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000,
		  120'b000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000,
		  120'b000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000,
		  120'b000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000,
		  120'b000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000,
		  120'b000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000,
		  120'b000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000,
		  120'b000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000,
		  120'b000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000,
		  120'b000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000,
		  120'b000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000,
		  120'b000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000,
		  120'b000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000,
		  120'b000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000,
		  120'b000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000,
		  120'b000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000000,
		  120'b000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000000,
		  120'b000000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000,
		  120'b000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000,
		  120'b000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000000,
		  120'b000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000,
		  120'b000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000,
		  120'b000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000,
		  120'b000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000,
		  120'b000000000000000000011111111111100000000000000000000000000000000000000000000000000000000001111111111110000000000000000000,
		  120'b000000000000000000011111111111110000000000000000000000000000000000000000000000000000000011111111111110000000000000000000,
		  120'b000000000000000000001111111111111100000000000000000000000000000000000000000000000000001111111111111100000000000000000000,
		  120'b000000000000000000000111111111111110000000000000000000000000000000000000000000000000011111111111111000000000000000000000,
		  120'b000000000000000000000011111111111111000000000000000000000000000000000000000000000000111111111111110000000000000000000000,
		  120'b000000000000000000000011111111111111100000000000000000000000000000000000000000000001111111111111110000000000000000000000,
		  120'b000000000000000000000001111111111111111000000000000000000000000000000000000000000111111111111111100000000000000000000000,
		  120'b000000000000000000000000111111111111111110000000000000000000000000000000000000011111111111111111000000000000000000000000,
		  120'b000000000000000000000000011111111111111111100000000000000000000000000000000001111111111111111110000000000000000000000000,
		  120'b000000000000000000000000001111111111111111111000000000000000000000000000000111111111111111111100000000000000000000000000,
		  120'b000000000000000000000000000011111111111111111111000000000000000000000000111111111111111111110000000000000000000000000000,
		  120'b000000000000000000000000000001111111111111111111111000000000000000000111111111111111111111100000000000000000000000000000,
		  120'b000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000,
		  120'b000000000000000000000000000000011111111111111111111111111111111111111111111111111111111110000000000000000000000000000000,
		  120'b000000000000000000000000000000000111111111111111111111111111111111111111111111111111111000000000000000000000000000000000,
		  120'b000000000000000000000000000000000011111111111111111111111111111111111111111111111111110000000000000000000000000000000000,
		  120'b000000000000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000000000,
		  120'b000000000000000000000000000000000000001111111111111111111111111111111111111111111100000000000000000000000000000000000000,
		  120'b000000000000000000000000000000000000000011111111111111111111111111111111111111110000000000000000000000000000000000000000,
		  120'b000000000000000000000000000000000000000000011111111111111111111111111111111110000000000000000000000000000000000000000000,
		  120'b000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000,
		  120'b000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,

         // code x02
        
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
		  120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000,
		  120'b000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000,
		  120'b000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000,  
		  120'b000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000,
		  120'b000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000,
		  120'b000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000,
		  120'b000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000,  
		  120'b000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000,  
		  120'b000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000,  
		  120'b000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000,  
		  120'b000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000,  
		  120'b000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000,  
		  120'b000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000,  
		  120'b000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000,  
		  120'b000000000000000000111111111111100000000000000000000000000000000000000000000000000000000001111111111111000000000000000000,  
		  120'b000000000000000000011111111111110000000000000000000000000000000000000000000000000000000011111111111110000000000000000000,  
		  120'b000000000000000000001111111111111000000000000000000000000000000000000000000000000000000111111111111100000000000000000000,  
		  120'b000000000000000000000111111111111100000000000000000000000000000000000000000000000000001111111111111000000000000000000000,  
		  120'b000000000000000000000011111111111110000000000000000000000000000000000000000000000000011111111111110000000000000000000000,  
		  120'b000000000000000000000001111111111111000000000000000000000000000000000000000000000000111111111111100000000000000000000000,  
		  120'b000000000000000000000000111111111111100000000000000000000000000000000000000000000001111111111111000000000000000000000000,  
		  120'b000000000000000000000000011111111111110000000000000000000000000000000000000000000011111111111110000000000000000000000000,  
		  120'b000000000000000000000000001111111111111000000000000000000000000000000000000000000111111111111100000000000000000000000000,  
		  120'b000000000000000000000000000111111111111100000000000000000000000000000000000000001111111111111000000000000000000000000000,  
		  120'b000000000000000000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000000000000000,  
		  120'b000000000000000000000000000001111111111111000000000000000000000000000000000000111111111111100000000000000000000000000000,  
		  120'b000000000000000000000000000000111111111111100000000000000000000000000000000001111111111111000000000000000000000000000000,  
		  120'b000000000000000000000000000000011111111111110000000000000000000000000000000011111111111110000000000000000000000000000000,  
		  120'b000000000000000000000000000000001111111111111000000000000000000000000000000111111111111100000000000000000000000000000000,  
		  120'b000000000000000000000000000000000111111111111100000000000000000000000000001111111111111000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000011111111111110000000000000000000000000011111111111110000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000001111111111111000000000000000000000000111111111111100000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000111111111111100000000000000000000001111111111111000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000011111111111110000000000000000000011111111111110000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000001111111111111000000000000000000111111111111100000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000111111111111100000000000000001111111111111000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000011111111111110000000000000011111111111110000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000001111111111111000000000000111111111111100000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000111111111111100000000001111111111111000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000011111111111110000000011111111111110000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000001111111111111000000111111111111100000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000000111111111111100001111111111111000000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000000011111111111110011111111111110000000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000,
		  120'b000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000000011111111111110011111111111110000000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000000111111111111100001111111111111000000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000001111111111111000000111111111111100000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000011111111111110000000011111111111110000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000000111111111111100000000001111111111111000000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000001111111111111000000000000111111111111100000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000011111111111110000000000000011111111111110000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000000111111111111100000000000000001111111111111000000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000001111111111111000000000000000000111111111111100000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000011111111111110000000000000000000011111111111110000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000000111111111111100000000000000000000001111111111111000000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000001111111111111000000000000000000000000111111111111100000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000011111111111110000000000000000000000000011111111111110000000000000000000000000000000000,  
		  120'b000000000000000000000000000000000111111111111100000000000000000000000000001111111111111000000000000000000000000000000000,  
		  120'b000000000000000000000000000000001111111111111000000000000000000000000000000111111111111100000000000000000000000000000000,  
		  120'b000000000000000000000000000000011111111111110000000000000000000000000000000011111111111110000000000000000000000000000000,  
		  120'b000000000000000000000000000000111111111111100000000000000000000000000000000001111111111111000000000000000000000000000000,  
		  120'b000000000000000000000000000001111111111111000000000000000000000000000000000000011111111111110000000000000000000000000000,  
		  120'b000000000000000000000000000011111111111110000000000000000000000000000000000000011111111111110000000000000000000000000000,  
		  120'b000000000000000000000000000111111111111100000000000000000000000000000000000000001111111111111000000000000000000000000000,  
		  120'b000000000000000000000000001111111111111000000000000000000000000000000000000000000111111111111100000000000000000000000000,  
		  120'b000000000000000000000000011111111111110000000000000000000000000000000000000000000011111111111110000000000000000000000000,  
		  120'b000000000000000000000000111111111111100000000000000000000000000000000000000000000001111111111111000000000000000000000000,  
		  120'b000000000000000000000001111111111111000000000000000000000000000000000000000000000000111111111111100000000000000000000000,  
		  120'b000000000000000000000011111111111110000000000000000000000000000000000000000000000000011111111111110000000000000000000000,  
		  120'b000000000000000000000111111111111100000000000000000000000000000000000000000000000000001111111111111000000000000000000000,  
		  120'b000000000000000000001111111111111000000000000000000000000000000000000000000000000000000111111111111100000000000000000000,  
		  120'b000000000000000000011111111111110000000000000000000000000000000000000000000000000000000011111111111110000000000000000000,  
		  120'b000000000000000000111111111111100000000000000000000000000000000000000000000000000000000001111111111111000000000000000000,  
		  120'b000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000,  
		  120'b000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000,  
		  120'b000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000,  
		  120'b000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000,  
		  120'b000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000,  
		  120'b000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000,  
		  120'b000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000,  
		  120'b000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000,  
		  120'b000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000,
		  120'b000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000,
		  120'b000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000,
		  120'b000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000,
		  120'b000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000,  
		  120'b000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 // 0
        };

	assign data = ROM[addr];

endmodule  
