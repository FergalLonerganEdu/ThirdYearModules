module lookuptable_rom_5 ( input [4:0]	addr,
						output [35:0]	data
					 );
				
	// ROM definition				
	parameter [0:27][35:0] ROM = {
	36'b010000011010100101010010011010100101,
	36'b010001011010100100011001011010100100,
	36'b010100101000000001010100101010000001, //p23
	36'b010001101000000001010001101010000001,
	36'b010000101000010001010000101010010001,
	36'b010000101000000101010000101010000101,
	36'b010000101001000001010010101001000001,
	36'b010110101001000001010110101001100001, //p23 part 2
	36'b010010101001000101010010101001100101,
	36'b010010101001010001010010101001011001,
	36'b000100011000000000100100011000000000, //p24
	36'b000100001000000100100100001000000100,
	36'b100101011000000000100101011000000010, //p26
	36'b100100011001000000100100011001000010,
	36'b100100011000010000100100011000010010,
	36'b100100011000000100100100011000000110,
	36'b100100011000000001100110011000000001,
	36'b100110011001000001100110011001100001, //p26 part 2
	36'b100110011000000101100110011000100101,
	36'b100110011000010001100110011000011001,
	36'b100101001000000100100101001000000110, //p28
	36'b100100011000000100100100011000000110,
	36'b100100001001000100100100001001000110,
	36'b100100001000010100100100001000010110,
	36'b100100001000000101100100001000100101,
	36'b100100011000100101100110011000100101, //p28 part 2
	36'b100100001001100101100110001001100101,
	36'b100101001000100101100101101000100101
};


assign data = ROM[addr];

endmodule  
