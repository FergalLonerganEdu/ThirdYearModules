module conor_rom ( input [11:0]	addr,
						output [23:0]	data
					 );

	parameter ADDR_WIDTH = 12;
   parameter DATA_WIDTH =  24;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2499][23:0] ROM = {
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfffffd,
		24'hfcfbff,
		24'hfffeff,
		24'hf7f9f4,
		24'hbabbb3,
		24'hb7b8b3,
		24'hbcbbb6,
		24'ha19f90,
		24'h9b9c8e,
		24'h9d9e90,
		24'h9b9b91,
		24'h8e8e86,
		24'h94938e,
		24'h81827d,
		24'h696a65,
		24'h686964,
		24'h6f6f6d,
		24'h747472,
		24'h6e6e6c,
		24'h6a6a6a,
		24'h666465,
		24'h6f6d6e,
		24'h868487,
		24'h686669,
		24'h64605f,
		24'h686860,
		24'h70716b,
		24'haaabb0,
		24'hfeffff,
		24'hfffffd,
		24'hfffffb,
		24'hfefcff,
		24'hffffff,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfdfcfa,
		24'hfffeff,
		24'hf9f8fd,
		24'hc2c4bf,
		24'hb4b5af,
		24'ha3a49f,
		24'ha2a19c,
		24'h959384,
		24'h8d8e7e,
		24'h9c9d8f,
		24'h919187,
		24'h77776f,
		24'h6d6c67,
		24'h61625c,
		24'h5c5d57,
		24'h5d5e58,
		24'h696a65,
		24'h63645f,
		24'h565752,
		24'h52534e,
		24'h555553,
		24'h626260,
		24'h777674,
		24'h5f5e5c,
		24'h535250,
		24'h52534e,
		24'h4f514e,
		24'h626367,
		24'hd0d1d5,
		24'hfeffff,
		24'hfefefe,
		24'hfefcff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfffffd,
		24'hfffeff,
		24'hd7d6db,
		24'ha0a29d,
		24'h969791,
		24'h91928d,
		24'h989792,
		24'h99978a,
		24'h989989,
		24'ha0a193,
		24'h84847a,
		24'h6b6b63,
		24'h5e5d58,
		24'h5c5d57,
		24'h63645e,
		24'h60615b,
		24'h5d6059,
		24'h575a53,
		24'h4f504a,
		24'h4d4e48,
		24'h4d4e49,
		24'h565752,
		24'h676863,
		24'h5f605b,
		24'h595856,
		24'h4e4e50,
		24'h48494d,
		24'h515254,
		24'h67686a,
		24'hc7c8cc,
		24'hfeffff,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfffffd,
		24'hecebf1,
		24'haeadb2,
		24'ha3a5a0,
		24'h888983,
		24'h888886,
		24'h8f8e89,
		24'h929083,
		24'ha8a99b,
		24'h96968a,
		24'h6f6f65,
		24'h66665e,
		24'h605f5a,
		24'h61625c,
		24'h61625c,
		24'h5a5b53,
		24'h555752,
		24'h545651,
		24'h555752,
		24'h555651,
		24'h4f504b,
		24'h50514c,
		24'h5e5f5a,
		24'h676863,
		24'h666664,
		24'h515056,
		24'h55545a,
		24'h474946,
		24'h3f4140,
		24'h67686d,
		24'he7e8ed,
		24'hfdfffc,
		24'hffffff,
		24'hfefefe,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfffeff,
		24'hc6c5cb,
		24'h8c8b91,
		24'h929491,
		24'h878883,
		24'h838381,
		24'h908f8b,
		24'h9e9c90,
		24'ha0a094,
		24'h7f7f75,
		24'h616159,
		24'h62615c,
		24'h605f5a,
		24'h5f605a,
		24'h585953,
		24'h575852,
		24'h585858,
		24'h555555,
		24'h585858,
		24'h5d5d5d,
		24'h5b5b5b,
		24'h5a5a5a,
		24'h636260,
		24'h706f6d,
		24'h6b6a66,
		24'h605e63,
		24'h4d4b50,
		24'h51514f,
		24'h454543,
		24'h43434b,
		24'ha1a1a9,
		24'hfcffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfaf8f9,
		24'h9a999f,
		24'h86858b,
		24'h8b8d8a,
		24'h7d7e79,
		24'h7b7b7b,
		24'h8b8a86,
		24'ha09e92,
		24'h8e8e84,
		24'h707068,
		24'h61605b,
		24'h61605c,
		24'h605f5b,
		24'h62635e,
		24'h5b5c57,
		24'h5c5d57,
		24'h595959,
		24'h575556,
		24'h5c5a5b,
		24'h686667,
		24'h6b6a68,
		24'h6a6967,
		24'h6b6a68,
		24'h777372,
		24'h71706c,
		24'h676364,
		24'h565253,
		24'h575352,
		24'h575556,
		24'h46454b,
		24'h64646c,
		24'heff2f7,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hf6f4f5,
		24'h7c7b83,
		24'h8e8d93,
		24'h989a99,
		24'h7b7c77,
		24'h787878,
		24'h8d8c88,
		24'h9b998d,
		24'h7d7c77,
		24'h676661,
		24'h62615d,
		24'h5e5d5b,
		24'h605f5d,
		24'h61615f,
		24'h5f5f5d,
		24'h5d5e59,
		24'h5a5955,
		24'h5d5956,
		24'h635f5c,
		24'h73706b,
		24'h76736e,
		24'h73706b,
		24'h706d68,
		24'h737069,
		24'h726e6b,
		24'h6a655f,
		24'h5a554f,
		24'h4c4646,
		24'h5c575b,
		24'h545255,
		24'h4a494f,
		24'hb1b1bd,
		24'hfcfcfc,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hfefefe,
		24'hffffff,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hf5f3f6,
		24'h7a7981,
		24'ha6a5ad,
		24'hb8bab9,
		24'ha4a5a0,
		24'h828282,
		24'h8b8a88,
		24'h838175,
		24'h6e6d69,
		24'h61605c,
		24'h62615f,
		24'h5f5d5e,
		24'h636162,
		24'h626262,
		24'h666664,
		24'h656563,
		24'h636059,
		24'h64615a,
		24'h67645b,
		24'h79756c,
		24'h7c786f,
		24'h79756a,
		24'h736f64,
		24'h716d62,
		24'h716c69,
		24'h676358,
		24'h60594f,
		24'h4f4647,
		24'h4f494d,
		24'h545051,
		24'h4e4d53,
		24'h676676,
		24'hf8f8f8,
		24'hfcfcfc,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hf4f4fe,
		24'h89868f,
		24'ha09798,
		24'haba49a,
		24'h9e9a8f,
		24'h908f8d,
		24'h898788,
		24'h7e7b74,
		24'h706c69,
		24'h6b6764,
		24'h6a6663,
		24'h6d6966,
		24'h6e6966,
		24'h787370,
		24'h746f6c,
		24'h726c6c,
		24'h6f6b68,
		24'h6a6663,
		24'h726f6a,
		24'h7c7974,
		24'h807d76,
		24'h7d7a73,
		24'h757269,
		24'h747168,
		24'h767269,
		24'h6a655f,
		24'h595450,
		24'h514d44,
		24'h514d41,
		24'h555146,
		24'h504d48,
		24'h504b4f,
		24'hb4b1c6,
		24'hfffeff,
		24'hfffffb,
		24'hfffffa,
		24'hfcfcfe,
		24'hfffeff,
		24'hfdfdfd,
		24'hfffffa,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hdcdfe8,
		24'h827f8a,
		24'haca3a6,
		24'hbcb5ad,
		24'ha9a49e,
		24'ha29da1,
		24'h969197,
		24'h898481,
		24'h7f7a77,
		24'h7f7a77,
		24'h807b78,
		24'h847f7c,
		24'h847f7c,
		24'h837e7b,
		24'h7f7a77,
		24'h827d7a,
		24'h7e7a77,
		24'h726e6b,
		24'h74716c,
		24'h787570,
		24'h77746d,
		24'h75726b,
		24'h706d64,
		24'h6d6a61,
		24'h6c685f,
		24'h6c6761,
		24'h5f5a57,
		24'h504b47,
		24'h4e4a41,
		24'h555249,
		24'h4f4b48,
		24'h4d484c,
		24'h625f72,
		24'hf5f4fc,
		24'hfffffb,
		24'hfffffb,
		24'hffffff,
		24'hfdfcff,
		24'hffffff,
		24'hfffffa,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hfdfdfd,
		24'hb4b8c1,
		24'h82808b,
		24'hbbb5b7,
		24'he4ddd7,
		24'hd6cecb,
		24'hbab3ba,
		24'h9e96a1,
		24'h988f92,
		24'h938b89,
		24'h908886,
		24'h8f8785,
		24'h8d8885,
		24'h8e8986,
		24'h8b8682,
		24'h8b8682,
		24'h87827e,
		24'h837e7b,
		24'h6f6a67,
		24'h67625e,
		24'h645f5b,
		24'h5e5955,
		24'h5e5953,
		24'h5f5a54,
		24'h5e5953,
		24'h656156,
		24'h66615d,
		24'h5b5555,
		24'h4e4848,
		24'h4c4845,
		24'h54504d,
		24'h4d4948,
		24'h4a4647,
		24'h555361,
		24'hf4f3f9,
		24'hfefefc,
		24'hfefffa,
		24'hffffff,
		24'hfcfbff,
		24'hffffff,
		24'hfefffa,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hfbfbfb,
		24'h848b91,
		24'h737479,
		24'hbeb8b8,
		24'hfff8f0,
		24'he8e1db,
		24'hb9b2b9,
		24'h9d939e,
		24'h968b91,
		24'h908788,
		24'h908788,
		24'h948c8a,
		24'h8c8784,
		24'h86817e,
		24'h87827e,
		24'h8d8a85,
		24'h817e79,
		24'h6f6a67,
		24'h615c59,
		24'h595451,
		24'h57524e,
		24'h544f4b,
		24'h55504c,
		24'h595450,
		24'h5b5650,
		24'h58544b,
		24'h595450,
		24'h5e5858,
		24'h5a5559,
		24'h4e494d,
		24'h4a4647,
		24'h474344,
		24'h4e4a49,
		24'ha4a2ad,
		24'hfffeff,
		24'hfffffd,
		24'hfefefc,
		24'hfdfdff,
		24'hfefdff,
		24'hffffff,
		24'hfffffd,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfdfdfd,
		24'hfbfbfb,
		24'h8d9598,
		24'h7b7c80,
		24'hc7c3c0,
		24'hece5db,
		24'haeaaa1,
		24'h8a8589,
		24'h7e777e,
		24'h716869,
		24'h71686b,
		24'h777173,
		24'h827c7c,
		24'h857f7f,
		24'h87827f,
		24'h85827d,
		24'h7e7b76,
		24'h6e6b64,
		24'h615c59,
		24'h5e5956,
		24'h5f5a57,
		24'h635e5b,
		24'h635e5b,
		24'h615c58,
		24'h635e5a,
		24'h65605c,
		24'h5e5953,
		24'h514c48,
		24'h575352,
		24'h5c575b,
		24'h4b464c,
		24'h443f45,
		24'h454044,
		24'h504c4d,
		24'hb0afb5,
		24'hfafafc,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfdfdff,
		24'hfcfcfc,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hfbfbfb,
		24'h889196,
		24'h797c81,
		24'hbdb9b8,
		24'hbbb7ac,
		24'h7f7c75,
		24'h727073,
		24'h6b696e,
		24'h635f5e,
		24'h636166,
		24'h6e696f,
		24'h716c70,
		24'h767273,
		24'h7a7675,
		24'h76726f,
		24'h67645f,
		24'h66615d,
		24'h696562,
		24'h686461,
		24'h66625f,
		24'h66625f,
		24'h615d5a,
		24'h5c5855,
		24'h605c59,
		24'h625e5b,
		24'h686560,
		24'h514e49,
		24'h524f4a,
		24'h555150,
		24'h49444a,
		24'h464148,
		24'h433e44,
		24'h454344,
		24'ha1a1a3,
		24'hffffff,
		24'hffffff,
		24'hfdfdfd,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hfcfcfc,
		24'h9ca4af,
		24'h828491,
		24'h99979c,
		24'h908d88,
		24'h777873,
		24'h77787d,
		24'h787880,
		24'h777777,
		24'h67676f,
		24'h6c6d72,
		24'h6d6c71,
		24'h686669,
		24'h595758,
		24'h5d5958,
		24'h57524f,
		24'h66615d,
		24'h6f6e6a,
		24'h686763,
		24'h656460,
		24'h63625e,
		24'h575652,
		24'h53524e,
		24'h5c5b59,
		24'h5c5b59,
		24'h64605f,
		24'h5a5752,
		24'h605d54,
		24'h5e5b56,
		24'h4d494a,
		24'h454047,
		24'h3b383f,
		24'h424043,
		24'ha4a4a2,
		24'hffffff,
		24'hffffff,
		24'hfcfcfe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hfdfdfd,
		24'ha3a8bb,
		24'h737488,
		24'h716e79,
		24'h81807e,
		24'h848484,
		24'h797c85,
		24'h80838c,
		24'h737478,
		24'h686b74,
		24'h676a71,
		24'h717277,
		24'h76757a,
		24'h646265,
		24'h736f6e,
		24'h66615e,
		24'h625d5a,
		24'h686763,
		24'h61605c,
		24'h666561,
		24'h6c6b67,
		24'h5f5e5c,
		24'h5e5d5b,
		24'h6a6967,
		24'h646361,
		24'h6b6768,
		24'h66635e,
		24'h69675b,
		24'h636057,
		24'h514d4c,
		24'h444148,
		24'h3c3940,
		24'h4b494e,
		24'hc7c8c3,
		24'hfdfdfb,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hfefefe,
		24'hfefeff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hbdbdc7,
		24'h605f6f,
		24'h615f6d,
		24'h747476,
		24'h767674,
		24'h7a7b7f,
		24'h7f7f89,
		24'h686b74,
		24'h61646b,
		24'h686b72,
		24'h727378,
		24'h7d7b80,
		24'h8e898d,
		24'h958f91,
		24'h807778,
		24'h5d5352,
		24'h5f5b58,
		24'h676360,
		24'h656460,
		24'h63625e,
		24'h696864,
		24'h6c6b67,
		24'h6e6b66,
		24'h706d68,
		24'h726d67,
		24'h67625c,
		24'h6f6764,
		24'h716966,
		24'h5a5250,
		24'h433f3c,
		24'h3c3b39,
		24'h5b5b59,
		24'hf8f8f8,
		24'hfcfcfc,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hf4f5fa,
		24'h777686,
		24'h605d70,
		24'h7b7984,
		24'h929196,
		24'h8a8991,
		24'h898991,
		24'h77787c,
		24'h6a6b70,
		24'h717277,
		24'h747378,
		24'h7e797d,
		24'ha59fa1,
		24'h9c9492,
		24'h847a79,
		24'h695e5c,
		24'h5c5753,
		24'h635e5a,
		24'h65625d,
		24'h67645f,
		24'h6c6964,
		24'h6e6b66,
		24'h6e6965,
		24'h6e6965,
		24'h726b63,
		24'h766f67,
		24'h79706b,
		24'h6e6462,
		24'h5a524f,
		24'h413d3a,
		24'h42413d,
		24'h91918f,
		24'hfcfcfc,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfafbfd,
		24'h72717f,
		24'h5f5b72,
		24'h9895a6,
		24'hb2b0bb,
		24'ha2a1a9,
		24'h97969b,
		24'h83847f,
		24'h7b797c,
		24'h79777a,
		24'h827e7f,
		24'h8c8686,
		24'hb4acaa,
		24'ha69b99,
		24'h867875,
		24'h736562,
		24'h605951,
		24'h625b55,
		24'h615c56,
		24'h645f59,
		24'h68635d,
		24'h6d6862,
		24'h746c69,
		24'h78706d,
		24'h7a7168,
		24'h7d746d,
		24'h7c736c,
		24'h706762,
		24'h5b5350,
		24'h3e3935,
		24'h56524f,
		24'hd4d3cf,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hf9f9fb,
		24'h7b7b87,
		24'h706f7f,
		24'h9c9ca4,
		24'hbababc,
		24'hb1afb4,
		24'ha19fa0,
		24'h9b9893,
		24'h8e8888,
		24'h958f8f,
		24'h9f9795,
		24'ha79d9b,
		24'hc4b9b5,
		24'hbcaeab,
		24'h857671,
		24'h786964,
		24'h6e645b,
		24'h6b6259,
		24'h706760,
		24'h756e66,
		24'h777068,
		24'h7a716a,
		24'h7f7671,
		24'h827773,
		24'h83796f,
		24'h7c7269,
		24'h7a7067,
		24'h726962,
		24'h58514b,
		24'h48433f,
		24'h827e7b,
		24'hfdf9f6,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hf9f9fb,
		24'h9c9ca6,
		24'h7d7d85,
		24'hd3d5d0,
		24'hc8cabf,
		24'hb1b0ab,
		24'ha8a2a2,
		24'h978f8d,
		24'ha79f9d,
		24'hbeb4b3,
		24'hbdb3b1,
		24'hc6bbb9,
		24'headcd9,
		24'hccbdb8,
		24'h877571,
		24'h786760,
		24'h71645c,
		24'h6b6158,
		24'h6e655c,
		24'h786f66,
		24'h7d746b,
		24'h80776e,
		24'h837970,
		24'h84776f,
		24'h83766d,
		24'h80736a,
		24'h7a7067,
		24'h6e675f,
		24'h524d47,
		24'h5a5752,
		24'hb8b4b1,
		24'hfffefd,
		24'hfefefe,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hedeef3,
		24'ha5a6a8,
		24'hd0d3c8,
		24'hd8dacc,
		24'hbdbab3,
		24'hb3aaad,
		24'hb7acb0,
		24'hafa5a4,
		24'hb2a6a6,
		24'hb1a6a4,
		24'hd4c6c5,
		24'hf8e9e6,
		24'hbdaba9,
		24'h8d7b77,
		24'h7a6864,
		24'h776966,
		24'h6c615d,
		24'h6b605a,
		24'h736a63,
		24'h7c736a,
		24'h83796f,
		24'h867c72,
		24'h877a71,
		24'h82746b,
		24'h80736b,
		24'h746b64,
		24'h6c655f,
		24'h524f4a,
		24'h5a5653,
		24'hd0cfcd,
		24'hfffffd,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfcfdf8,
		24'hfeffff,
		24'hf3f4f9,
		24'ha6a8a3,
		24'hcbccc6,
		24'hc9c5c4,
		24'hc1b6bc,
		24'hbbafb3,
		24'hb9adaf,
		24'ha4989a,
		24'ha99b9b,
		24'hc5b7b7,
		24'hd0c0c0,
		24'ha08e8e,
		24'h8e7c7a,
		24'h7b6967,
		24'h746666,
		24'h6e6361,
		24'h6f6460,
		24'h756c65,
		24'h7c736a,
		24'h80766c,
		24'h80766a,
		24'h817567,
		24'h81726b,
		24'h786e65,
		24'h6d665e,
		24'h6a655f,
		24'h51504c,
		24'h4b4a48,
		24'hd6d4d5,
		24'hfffdfe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfffff6,
		24'hfbfcff,
		24'hfefeff,
		24'ha0a1a6,
		24'hb5b4b9,
		24'hc0bbc2,
		24'hc2b7bf,
		24'hc2b3b6,
		24'hb5a9ab,
		24'hab9fa1,
		24'haa9b9e,
		24'ha09292,
		24'h948485,
		24'h8d7d7e,
		24'h837171,
		24'h766464,
		24'h695a5d,
		24'h6a5e5e,
		24'h6f6563,
		24'h766d68,
		24'h7a7168,
		24'h7b7366,
		24'h7e7566,
		24'h847868,
		24'h7d7068,
		24'h736960,
		24'h6e675f,
		24'h686560,
		24'h4d4e49,
		24'h454543,
		24'hdbdbdb,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfdfffe,
		24'hfeffff,
		24'hd5d9dc,
		24'h9a9da4,
		24'hb8b7bd,
		24'hbebcbd,
		24'hb8b5b0,
		24'hb6acad,
		24'hb1a5a5,
		24'hbeb0af,
		24'had9e9b,
		24'h998a87,
		24'h8d7e7b,
		24'h7e6e6e,
		24'h746666,
		24'h695f5d,
		24'h695f5d,
		24'h716863,
		24'h797069,
		24'h796f66,
		24'h796f65,
		24'h7d7367,
		24'h7d7367,
		24'h787065,
		24'h71685f,
		24'h6d645d,
		24'h6b6360,
		24'h504b48,
		24'h525051,
		24'hefeff1,
		24'hfeffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfbfdfc,
		24'hfeffff,
		24'hf9fdff,
		24'hdfe0e5,
		24'hc2c1c7,
		24'hc1c0be,
		24'hbcb9b4,
		24'hb6b1ae,
		24'hbdb5b3,
		24'hc9bfbd,
		24'hc6bbb7,
		24'hb6a8a5,
		24'h948685,
		24'h7d7270,
		24'h776b6b,
		24'h736866,
		24'h706561,
		24'h716662,
		24'h736862,
		24'h736960,
		24'h746a60,
		24'h776d61,
		24'h776d61,
		24'h756d62,
		24'h6e655c,
		24'h716861,
		24'h635b58,
		24'h4d4845,
		24'h6b696a,
		24'hfefeff,
		24'hfeffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfdfdff,
		24'hfdfffe,
		24'hfeffff,
		24'hfafbfd,
		24'hfeffff,
		24'hcccbd0,
		24'hb8b8b8,
		24'hc2c1bc,
		24'hbebbb6,
		24'hbcb9b2,
		24'hb4ada7,
		24'hbab1ac,
		24'hb8ada9,
		24'h958a88,
		24'h827676,
		24'h7e7274,
		24'h827370,
		24'h7b6c69,
		24'h71645e,
		24'h6c5f59,
		24'h6f625a,
		24'h746a60,
		24'h7a7066,
		24'h7b7165,
		24'h6e675d,
		24'h6f685e,
		24'h6e675f,
		24'h5d5552,
		24'h4e4946,
		24'h939290,
		24'hfcfcfc,
		24'hfeffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfafcf9,
		24'hfdfffe,
		24'hfdfeff,
		24'hcfced3,
		24'hc3c3c1,
		24'hc5c6c0,
		24'hc8c5bc,
		24'hb3b0a7,
		24'h99928c,
		24'ha19893,
		24'haa9f9d,
		24'h968888,
		24'h887a7a,
		24'h807174,
		24'h796765,
		24'h746260,
		24'h6b5c57,
		24'h6b5c55,
		24'h72655d,
		24'h776d63,
		24'h796f65,
		24'h776f62,
		24'h6e675d,
		24'h6f6860,
		24'h645d55,
		24'h544c49,
		24'h4e4946,
		24'hcac9c7,
		24'hfefefe,
		24'hfeffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hfefefc,
		24'hffffff,
		24'hfefeff,
		24'hdedee0,
		24'haaacab,
		24'hbfc2bb,
		24'hcac8bc,
		24'ha5a198,
		24'h887f7a,
		24'h8d827e,
		24'h938383,
		24'h8a7779,
		24'h837072,
		24'h7e6b6d,
		24'h7c6a66,
		24'h776561,
		24'h71625d,
		24'h75665f,
		24'h7b6e66,
		24'h7c7268,
		24'h796f65,
		24'h766e63,
		24'h69655a,
		24'h67635a,
		24'h635c56,
		24'h4e4945,
		24'h56514e,
		24'heeedeb,
		24'hffffff,
		24'hfdfffe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfdfeff,
		24'hfdfdfd,
		24'hfffffb,
		24'hfbfaf8,
		24'hffffff,
		24'hf7f7f9,
		24'h9b9d9c,
		24'hb0b5af,
		24'hc0c0b4,
		24'ha3a097,
		24'h968f89,
		24'ha29795,
		24'ha49494,
		24'h998787,
		24'h8a7878,
		24'h837171,
		24'h7c6d68,
		24'h786964,
		24'h756860,
		24'h786b63,
		24'h7b6e66,
		24'h796f65,
		24'h766c62,
		24'h73695f,
		24'h656158,
		24'h5e5a51,
		24'h5b5650,
		24'h544f4b,
		24'h827e7b,
		24'hfffffd,
		24'hfefefe,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfeffff,
		24'hffffff,
		24'hfffefa,
		24'hfffffb,
		24'hfffeff,
		24'hffffff,
		24'hd3d7d6,
		24'h949993,
		24'ha8aea2,
		24'ha3a69d,
		24'h999893,
		24'h9f9a96,
		24'h9d9391,
		24'h928483,
		24'h7f716e,
		24'h746761,
		24'h736960,
		24'h746a61,
		24'h7a7067,
		24'h7e746b,
		24'h7c7268,
		24'h7a7066,
		24'h756b61,
		24'h6e645a,
		24'h625f56,
		24'h57534a,
		24'h524d47,
		24'h5c5753,
		24'h979390,
		24'hfffffd,
		24'hfffffd,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfdfeff,
		24'hfefefe,
		24'hfffefa,
		24'hfffffb,
		24'hfffdfe,
		24'hfefeff,
		24'hf6faf9,
		24'h747b74,
		24'h879387,
		24'ha5ada2,
		24'ha6a9a2,
		24'ha6a5a1,
		24'ha7a29e,
		24'h9f9892,
		24'h8e857e,
		24'h837a71,
		24'h7b7269,
		24'h7d746b,
		24'h827970,
		24'h80776e,
		24'h7a7066,
		24'h776d63,
		24'h72685e,
		24'h695f55,
		24'h58554c,
		24'h57544d,
		24'h5c5751,
		24'h625d59,
		24'h6b6764,
		24'hd6d5d3,
		24'hfffffd,
		24'hfdfdfd,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hfdfdfd,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfbffff,
		24'hfcffff,
		24'hfefeff,
		24'hffffff,
		24'hfcfcfe,
		24'hffffff,
		24'hfafeff,
		24'hcdd1d2,
		24'h737f7f,
		24'h93989b,
		24'hb2b0b1,
		24'hbcb4b1,
		24'hc4bbb2,
		24'hc9c1b6,
		24'hb2a7a1,
		24'h958a88,
		24'h878378,
		24'h858178,
		24'h7e7a71,
		24'h77736a,
		24'h747067,
		24'h716a62,
		24'h665f57,
		24'h5b544c,
		24'h534f4c,
		24'h54514c,
		24'h68655e,
		24'h6a6762,
		24'h615f60,
		24'ha7a6ac,
		24'hfeffff,
		24'hfcffff,
		24'hfefffa,
		24'hfdfef9,
		24'hffffff,
		24'hfffeff,
		24'hfcfbff,
		24'hffffff,
		24'hfdfdfd,
		24'hfefffd,
		24'hffffff,
		24'hfdfdfd,
		24'hfdfdfd,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hfdfdfd,
		24'hfefefe,
		24'hfffffd,
		24'hfffffd,
		24'hfefaf9,
		24'hfffefd,
		24'hfffefd,
		24'hfcf8f7,
		24'hfffffd,
		24'hfefefc,
		24'hafb3b4,
		24'h6b6f72,
		24'h999d9e,
		24'hb7bcb6,
		24'hb1b4a9,
		24'hacaca0,
		24'ha39a93,
		24'h908281,
		24'h848178,
		24'h7d7a71,
		24'h77736a,
		24'h716d64,
		24'h69645e,
		24'h5d5852,
		24'h544f49,
		24'h514c46,
		24'h544f4b,
		24'h646057,
		24'h6d6960,
		24'h706b65,
		24'h5f5b5c,
		24'h7d7a81,
		24'heff0f5,
		24'hfcffff,
		24'hfffffd,
		24'hfffffd,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfcfcfe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfdfdfb,
		24'hfffffd,
		24'hfffffd,
		24'hfffdfc,
		24'hfffefd,
		24'hfffffd,
		24'hfffffd,
		24'hfffffd,
		24'hf9fafc,
		24'h8b8f92,
		24'h7b8083,
		24'h8b918f,
		24'h868b84,
		24'h7b7c74,
		24'h807d76,
		24'h7e7975,
		24'h75726b,
		24'h6d6a63,
		24'h65625b,
		24'h615e57,
		24'h5a5750,
		24'h534e48,
		24'h544f49,
		24'h59544e,
		24'h676056,
		24'h716b5f,
		24'h767064,
		24'h777068,
		24'h696363,
		24'h5e595f,
		24'h8c8b93,
		24'hf7f8fd,
		24'hfffdff,
		24'hfcfafb,
		24'hfffffd,
		24'hfcfbf7,
		24'hfffffb,
		24'hfffffd,
		24'hfffeff,
		24'hfcfafd,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfcfffd,
		24'hfcfffd,
		24'hfefffd,
		24'hfdfffc,
		24'hfcfefb,
		24'hfdfffc,
		24'hfbfffc,
		24'hfbfffc,
		24'hfbfffe,
		24'hf1f5f8,
		24'hadaeb3,
		24'haeacaf,
		24'h85817e,
		24'h66635c,
		24'h5a5b53,
		24'h5c635b,
		24'h5f5c57,
		24'h595651,
		24'h55524d,
		24'h54514c,
		24'h54514c,
		24'h595651,
		24'h635e5a,
		24'h6a6561,
		24'h716b5d,
		24'h797262,
		24'h7a7363,
		24'h797268,
		24'h6e6566,
		24'h5d585e,
		24'h4f4c55,
		24'h95949c,
		24'hfbf9fe,
		24'hfffeff,
		24'hfffffb,
		24'hfefff9,
		24'hfefff7,
		24'hfefff9,
		24'hfffffd,
		24'hfffeff,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hfefefe,
		24'hfdfdfd,
		24'hffffff,
		24'hfbfcfe,
		24'hfeffff,
		24'hfeffff,
		24'hfdfeff,
		24'hfeffff,
		24'hfdfeff,
		24'hffffff,
		24'hfefefe,
		24'hfeffff,
		24'hdedfe3,
		24'hd6d2d3,
		24'hc3bbb8,
		24'ha59c97,
		24'h79766f,
		24'h6f716c,
		24'h6e6a67,
		24'h65615e,
		24'h615d5a,
		24'h63605b,
		24'h66635e,
		24'h6c6763,
		24'h726d69,
		24'h76716b,
		24'h7c7467,
		24'h7f7868,
		24'h7d7666,
		24'h776e65,
		24'h766e6c,
		24'h6e676e,
		24'h5b555f,
		24'h454249,
		24'h878588,
		24'hf2f0f3,
		24'hffffff,
		24'hfefffd,
		24'hfcfef9,
		24'hfefffa,
		24'hfdfcf8,
		24'hfefdf9,
		24'hffffff,
		24'hfefefe,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfdfdfd,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hfffdff,
		24'hfffdff,
		24'hfffdff,
		24'hfdfbfe,
		24'hfffdff,
		24'hfffeff,
		24'hfffcff,
		24'hfffdff,
		24'hfffdff,
		24'hfdfffe,
		24'hf3fcf7,
		24'hd7ded6,
		24'hd2d0c4,
		24'hc4bbb2,
		24'haca19d,
		24'h938b89,
		24'h837f7c,
		24'h736e6b,
		24'h6c6763,
		24'h716c68,
		24'h736e6a,
		24'h726d67,
		24'h76716b,
		24'h7a756f,
		24'h847c6f,
		24'h817a6a,
		24'h7d7666,
		24'h7c736a,
		24'h736b69,
		24'h625b62,
		24'h4f4c53,
		24'h444148,
		24'h454348,
		24'h78777d,
		24'hadadb9,
		24'hf8faff,
		24'hf9fbff,
		24'hfeffff,
		24'hffffff,
		24'hfffffb,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hfdfdfd,
		24'hffffff,
		24'hffffff,
		24'hfcfcfc,
		24'hfffffb,
		24'hfafcf7,
		24'hfbfffa,
		24'hfbfffb,
		24'hfbfffb,
		24'hfafff9,
		24'hfafcf7,
		24'hf1f2ed,
		24'heeeeec,
		24'hebf4ef,
		24'hc2d2c5,
		24'hddead8,
		24'hd8d9c7,
		24'hc5bcad,
		24'hb8aba5,
		24'h988e8d,
		24'h898481,
		24'h797470,
		24'h736e6a,
		24'h7a726f,
		24'h7b746e,
		24'h7c756f,
		24'h827b73,
		24'h878078,
		24'h868074,
		24'h877f72,
		24'h7e7669,
		24'h7b746a,
		24'h615957,
		24'h4d484e,
		24'h49464d,
		24'h47464c,
		24'h44434b,
		24'h414050,
		24'h494965,
		24'h707394,
		24'ha5a8c7,
		24'hf3f4ff,
		24'hfefeff,
		24'hfffffd,
		24'hfdfdfd,
		24'hffffff,
		24'hffffff,
		24'hfefefe,
		24'hffffff,
		24'hfefefe,
		24'hffffff,
		24'hffffff,
		24'hf9f9f9,
		24'hededed,
		24'hd1dfd2,
		24'hd5e5d8,
		24'he1f3e5,
		24'hdff4e5,
		24'hd3e8d9,
		24'hd0e2d4,
		24'haabaad,
		24'h616f62,
		24'h697871,
		24'hacc0b5,
		24'he5fae9,
		24'hf1fbe3,
		24'hded9c3,
		24'hc6baaa,
		24'hb4aba4,
		24'h9d9c9a,
		24'h918986,
		24'h88807d,
		24'h847c79,
		24'h847d77,
		24'h837c76,
		24'h877e77,
		24'h8b827b,
		24'h8c837a,
		24'h898278,
		24'h7b7569,
		24'h706a5e,
		24'h524b43,
		24'h4f4949,
		24'h4a454b,
		24'h49464d,
		24'h47464b,
		24'h4a4856,
		24'h434159,
		24'h3e3d65,
		24'h39396b,
		24'h414272,
		24'h78789a,
		24'h9c9ba9,
		24'hadadaf,
		24'hf5f5f5,
		24'hfafafa,
		24'hfefdfb,
		24'hffffff,
		24'hf9fafc,
		24'hfcffff,
		24'hfbffff,
		24'he0e8eb,
		24'hc1c9d4,
		24'hbcc3d6,
		24'hb3c1c2,
		24'hbccbc8,
		24'hc3d0c9,
		24'hbfccc5,
		24'hb6c1bd,
		24'ha7b0ad,
		24'h8e9890,
		24'h798378,
		24'hdcdadd,
		24'hfffffa,
		24'hffffef,
		24'hfffce3,
		24'he4dec6,
		24'hc6baaa,
		24'hbbaca7,
		24'had9d9e,
		24'h9d948d,
		24'h968d86,
		24'h948b84,
		24'h8f887e,
		24'h888276,
		24'h888478,
		24'h878377,
		24'h7b796a,
		24'h66665c,
		24'h535349,
		24'h474641,
		24'h474644,
		24'h48464b,
		24'h45424b,
		24'h46434e,
		24'h4a4654,
		24'h48465e,
		24'h4a485e,
		24'h49475c,
		24'h434254,
		24'h3f3e50,
		24'h413f54,
		24'h46445a,
		24'h49475f,
		24'h595762,
		24'h84828d,
		24'hfefefc,
		24'hffffff,
		24'hfeffff,
		24'hf4f8fb,
		24'hcbd0d3,
		24'hb8c0c3,
		24'hb3bcc5,
		24'habb2c2,
		24'ha9b4ba,
		24'ha4afb1,
		24'ha3adac,
		24'ha4aead,
		24'ha2aaad,
		24'h99a1a4,
		24'h929898,
		24'h8f9591,
		24'hc5c6be,
		24'he8e9db,
		24'hf9fbe5,
		24'hfbfbdf,
		24'hdeddc1,
		24'hbfbaa4,
		24'hada598,
		24'ha79c96,
		24'h9b9390,
		24'h928a87,
		24'h8a8581,
		24'h817c76,
		24'h737069,
		24'h69665d,
		24'h5d5d53,
		24'h505044,
		24'h4d4c4a,
		24'h464445,
		24'h464447,
		24'h49464d,
		24'h494651,
		24'h464251,
		24'h474354,
		24'h484357,
		24'h4a495b,
		24'h4a4959,
		24'h484755,
		24'h464652,
		24'h444450,
		24'h444351,
		24'h444353,
		24'h444355,
		24'h3f3f49,
		24'h4e4e58,
		24'hfefffb,
		24'hfafcfb,
		24'hdee1e6,
		24'hc3c6cd,
		24'hb2b7bd,
		24'habb2b8,
		24'ha3acb3,
		24'ha6aeb9,
		24'ha3abb6,
		24'ha4adb4,
		24'ha5acb2,
		24'h9fa6ac,
		24'h979ba4,
		24'h8d919a,
		24'h898c91,
		24'h878b8c,
		24'h7f8176,
		24'h828477,
		24'h8b8e7d,
		24'h929381,
		24'h8e8f7d,
		24'h868779,
		24'h77746b,
		24'h726f68,
		24'h6c6869,
		24'h626061,
		24'h5b595a,
		24'h575654,
		24'h50504e,
		24'h4c4d48,
		24'h4a4b46,
		24'h464843,
		24'h48474c,
		24'h48474c,
		24'h4b4a50,
		24'h4c4b53,
		24'h494752,
		24'h474552,
		24'h474553,
		24'h474553,
		24'h484852,
		24'h47474f,
		24'h47474f,
		24'h48494e,
		24'h494a4f,
		24'h494951,
		24'h484850,
		24'h484852,
		24'h494953,
		24'h4e4e58,
		24'hf8fdf7,
		24'hdadedf,
		24'hbabdc6,
		24'ha7abb6,
		24'ha3a7b2,
		24'ha4abb1,
		24'ha5acb2,
		24'ha6afb6,
		24'ha0a6b2,
		24'h9ea5ad,
		24'h989fa5,
		24'h8d9298,
		24'h82858e,
		24'h7e808c,
		24'h83838b,
		24'h848589,
		24'h848685,
		24'h747675,
		24'h6c6e6d,
		24'h656766,
		24'h5f6062,
		24'h5b5f60,
		24'h525659,
		24'h4f5356,
		24'h525358,
		24'h4f5055,
		24'h4d4e52,
		24'h4c4d51,
		24'h4b4f52,
		24'h494d50,
		24'h484c4d,
		24'h484c4d,
		24'h4c4c4e,
		24'h4b4b4d,
		24'h4b4b4d,
		24'h4a4a4c,
		24'h48474c,
		24'h48474c,
		24'h49484d,
		24'h48474c,
		24'h48494e,
		24'h48494e,
		24'h494a4e,
		24'h4a4b4f,
		24'h48494d,
		24'h45464a,
		24'h46474c,
		24'h4a4b50,
		24'h494951,
		24'h54545c,
		24'hd3d9d5,
		24'haeb3b6,
		24'h9fa3ae,
		24'h9a9dac,
		24'h9097a1,
		24'h92999f,
		24'h99a1a4,
		24'h98a0a3,
		24'h979ea8,
		24'h8c9399,
		24'h868b8f,
		24'h83888c,
		24'h80838a,
		24'h7e7e88,
		24'h7d7e83,
		24'h7d7e80,
		24'h77787d,
		24'h74777e,
		24'h767982,
		24'h727480,
		24'h676b76,
		24'h5d616c,
		24'h565d67,
		24'h4f5660,
		24'h4c4f56,
		24'h4e5158,
		24'h4d5057,
		24'h4d5057,
		24'h4d5258,
		24'h4b5054,
		24'h474c50,
		24'h454a4e,
		24'h4b4c50,
		24'h48494d,
		24'h48494d,
		24'h4a4b4d,
		24'h494a4c,
		24'h48494b,
		24'h494a4c,
		24'h48494b,
		24'h474a4f,
		24'h474a4f,
		24'h484b50,
		24'h484b50,
		24'h43464b,
		24'h3f4247,
		24'h414449,
		24'h46494e,
		24'h474a4f,
		24'h505358,
		24'hafb8b7,
		24'h99a0a6,
		24'h8c929e,
		24'h888e9c,
		24'h8e959f,
		24'h8d949a,
		24'h878f92,
		24'h8a9295,
		24'h858c94,
		24'h7a8285,
		24'h757a7d,
		24'h73787b,
		24'h74777e,
		24'h787b82,
		24'h7d7e83,
		24'h7c7d7f,
		24'h73777a,
		24'h707378,
		24'h6a6d72,
		24'h666b71,
		24'h656a70,
		24'h61666c,
		24'h5f666c,
		24'h545c5f,
		24'h4f545a,
		24'h50555b,
		24'h4d5258,
		24'h4b5056,
		24'h4b5056,
		24'h4d5057,
		24'h4b5056,
		24'h4a4f55,
		24'h4c4f58,
		24'h494c53,
		24'h4a4d54,
		24'h4c4f56,
		24'h494c53,
		24'h484b52,
		24'h484b50,
		24'h494c51,
		24'h484b50,
		24'h474a4f,
		24'h484b52,
		24'h494c53,
		24'h474a51,
		24'h44474e,
		24'h45484d,
		24'h484b50,
		24'h494d50,
		24'h505457,
		24'h97a1a3,
		24'h879097,
		24'h848c97,
		24'h808692,
		24'h818890,
		24'h7f878a,
		24'h7c8487,
		24'h7d848a,
		24'h787f89,
		24'h737a80,
		24'h70787b,
		24'h6e7377,
		24'h6b6f78,
		24'h6f727b,
		24'h72757c,
		24'h717277,
		24'h6f7277,
		24'h707477,
		24'h6f7376,
		24'h6c7073,
		24'h6d7174,
		24'h686e6e,
		24'h656b6b,
		24'h595f5f,
		24'h54575c,
		24'h52555a,
		24'h515459,
		24'h52555a,
		24'h52555a,
		24'h53565b,
		24'h53565b,
		24'h52555a,
		24'h4f5458,
		24'h4c5155,
		24'h4b5054,
		24'h4a4f53,
		24'h484d51,
		24'h484d51,
		24'h4b5054,
		24'h4b5054,
		24'h4b4f52,
		24'h4a4e51,
		24'h4a4d52,
		24'h4a4d54,
		24'h494c53,
		24'h474a4f,
		24'h484c4f,
		24'h4a4e51,
		24'h4c5053,
		24'h565a5d,
		24'h899299,
		24'h7b848d,
		24'h7d8590,
		24'h7a838c,
		24'h7d848a,
		24'h7a8285,
		24'h788083,
		24'h7a8189,
		24'h767e89,
		24'h697078,
		24'h666d73,
		24'h6c7079,
		24'h696d78,
		24'h656774,
		24'h656773,
		24'h676a71,
		24'h666972,
		24'h6a6d74,
		24'h717479,
		24'h6e7275,
		24'h727679,
		24'h707477,
		24'h6b6f72,
		24'h64686b,
		24'h606467,
		24'h595d60,
		24'h575b5e,
		24'h5a5b5f,
		24'h58595d,
		24'h57585c,
		24'h58595d,
		24'h595a5f,
		24'h575d59,
		24'h535955,
		24'h4f5551,
		24'h4c524e,
		24'h4a504c,
		24'h4c524e,
		24'h4c524e,
		24'h4a504c,
		24'h4a4e4d,
		24'h4a4e4f,
		24'h494d50,
		24'h484b50,
		24'h46494e,
		24'h464a4d,
		24'h494d4e,
		24'h4c504f,
		24'h4a5050,
		24'h535959,
		24'h7f8289,
		24'h747881,
		24'h818590,
		24'h81858e,
		24'h7b8084,
		24'h7a7f82,
		24'h797e82,
		24'h777c82,
		24'h757984,
		24'h6c7079,
		24'h6b6e77,
		24'h6a6d76,
		24'h666972,
		24'h666670,
		24'h65656f,
		24'h696973,
		24'h696a6f,
		24'h6d6e73,
		24'h717277,
		24'h707175,
		24'h6e6f73,
		24'h6d6e72,
		24'h6b6c6e,
		24'h696a6c,
		24'h636768,
		24'h5e6265,
		24'h5a5e61,
		24'h595c61,
		24'h585b60,
		24'h565a5d,
		24'h565a5d,
		24'h595d5e,
		24'h5c5e5d,
		24'h585a59,
		24'h525655,
		24'h505455,
		24'h4d5152,
		24'h4d5152,
		24'h4c5053,
		24'h4a4e51,
		24'h494d4e,
		24'h4a4e4f,
		24'h484c4d,
		24'h484c4d,
		24'h4a4e4f,
		24'h4a4e4d,
		24'h4a4e4d,
		24'h4b4f4e,
		24'h4a4e4d,
		24'h4b4f4e,
		24'h888b92,
		24'h7c8089,
		24'h878b96,
		24'h848891,
		24'h7e8387,
		24'h7e8386,
		24'h7f8488,
		24'h7d848a,
		24'h7d8285,
		24'h787d80,
		24'h777b7e,
		24'h727679,
		24'h6f7376,
		24'h737476,
		24'h737476,
		24'h727375,
		24'h74757a,
		24'h76777c,
		24'h77787d,
		24'h737478,
		24'h707175,
		24'h6f7074,
		24'h6e6f71,
		24'h6d6e70,
		24'h696d6e,
		24'h6b6f72,
		24'h696d70,
		24'h65686d,
		24'h62656a,
		24'h616568,
		24'h616568,
		24'h5f6364,
		24'h626463,
		24'h5e605f,
		24'h5b5f5e,
		24'h595d5e,
		24'h585c5d,
		24'h575b5c,
		24'h575b5e,
		24'h54585b,
		24'h535758,
		24'h535758,
		24'h525657,
		24'h525657,
		24'h545859,
		24'h545857,
		24'h545857,
		24'h555958,
		24'h545857,
		24'h5c605f
	};

	assign data = ROM[addr];

endmodule  
