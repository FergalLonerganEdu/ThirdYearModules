module lookuptable_rom_4 ( input [4:0]	addr,
						output [35:0]	data
					 );

	// ROM definition				
	parameter [0:27][35:0] ROM = {
	36'b010001001000000000011001001000000000,
	36'b010000011000000000010000011000100000,
	36'b010000001000000100010000001010000100,
	36'b010000001000010000010000101000010000,
	36'b010000001001000000010000001001001000,
	36'b010000001000000001010000101000000001,
	36'b010110011000000000010110011000100000, //p20
	36'b010110001001000000010110001001100000,
	36'b010110001000000100010110001000000100,
	36'b010110001000000001010110001000100001,
	36'b010110001000010000010110101000010000,
	36'b010110101000010100010110101010010100, //p20 part 2
	36'b010110101000010001010110101010010001,
	36'b010110101001010000010110101001010010,
	36'b011001011000000000011001011000001000, //p21
	36'b011001001000010000011001001000011000,
	36'b011001001001000000011001001001001000,
	36'b011001001000000001001001001000001001,
	36'b011001001000000100011001001000100100,
	36'b011001001000100101011001001010100101, //p21 part 2
	36'b011001001001100100011001001001100110,
	36'b011001011000100100011001011010100100,
	36'b010100001010000100010100101010000100, //p22
	36'b010001001010000100010001101010000100,
	36'b010000001010010100010000101010010100,
	36'b010000001010000101010000101010000101,
	36'b010000011010000100010000011010100100,
	36'b010100011010100100010110011010100100  //p22 part 2
};


assign data = ROM[addr];

endmodule  
