module lookuptable_rom_2 ( input [4:0]	addr,
						output [35:0]	data
					 );
				
	// ROM definition				
	parameter [0:27][35:0] ROM = {
	36'b000110100100011001100110100100011001, //p8
	36'b000110100101011000000110100101011010,
	36'b010110100100011000010110100100011010,
	36'b010110010110001000010110010110001010, //p9
	36'b000110010110011000010110010110001010,
	36'b000110010110001001100110010110001001,
	36'b010110100101001000010110100101001010, //p10
	36'b000110100101011000000110100101011010,
	36'b000100000000000000000100001000000000,
	36'b010010010110000000010010010110000010, //p11
	36'b000110010110000000000110000010000010,
	36'b000010010110010000000010010110010010,
	36'b000010010110000100000010010110000110,
	36'b000010010110000001100010010110000001,
	36'b100010010110010001101010010110010001, //p11 part 2
	36'b100010010110000101101010010110000101,
	36'b100110010110000001100110010110001001,
	36'b100010010100010000101010010100010000, //p12
	36'b100010000101010000101010000101010000,
	36'b100010000100010100101010000100010100,
	36'b100010000100010001101010000100010001,
	36'b100110000100010000100110000100011000,
	36'b100110010100011000100110010110011000, //p12 part 2
	36'b100110000101011000100110100101011000,
	36'b100110000100011001100110100100011001,
	36'b001010010100000100101010010100000100, //p13
	36'b001010000100010100101010000100010100,
	36'b001010000101000100101010000101000100
};


assign data = ROM[addr];

endmodule  
