module lookuptable_rom_3 ( input [4:0]	addr,
						output [35:0]	data
					 );
				
	// ROM definition				
	parameter [0:27][35:0] ROM = {
	36'b001010000100000101101010000100000101,
	36'b011010000100000100011010000100000110,
	36'b011010010100000110011010010110000110, //p13 part 2
	36'b011010000101000110011010100101000110,
	36'b011010000100010110011010000110010110,
	36'b100010010100000001101010010100000001, //p14
	36'b100010000100010001101010000100010001,
	36'b100010000100000101101010000100000101,
	36'b100010000101000001101010000101000001,
	36'b100110000100000001100110000100001001,
	36'b100110010100001001100110010110001001, //p14 part 2
	36'b100110000101001001100110100101001001,
	36'b100110000100011001100110000110011001,
	36'b000110100101000000000110100101001000, //p15
	36'b010010100101000000010010100101000010,
	36'b000010100101010000100010100101010000,
	36'b000010100101000100001010100101000100,
	36'b000010100101000001100010100101000001,
	36'b100010100101010100101010100101010100, //p16
	36'b100010100101010001101010100101010001,
	36'b100110100101010000100110100101011000,
	36'b001010100101010100101010100101010100, //p17
	36'b001010100101000101101010100101000101,
	36'b011010100101000100011010100101000110,
	36'b100010100101010001101010100101010001, //p18
	36'b100010100101000101101010100101000101,
	36'b100110100101000001100110100101100001,
	36'b010100001000000000010110001000000000 //p19
};


assign data = ROM[addr];

endmodule  
