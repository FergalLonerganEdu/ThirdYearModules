module sprite_addr_rom (input [5:0] xcoord, ycoord,
								output logic [11:0] addr);

	logic [5:0] xcoord_reg;
	logic [5:0] ycoord_reg;
	parameter [0:49][0:49][11:0] ROM = {
		12'h000,
		12'h001,
		12'h002,
		12'h003,
		12'h004,
		12'h005,
		12'h006,
		12'h007,
		12'h008,
		12'h009,
		12'h00a,
		12'h00b,
		12'h00c,
		12'h00d,
		12'h00e,
		12'h00f,
		12'h010,
		12'h011,
		12'h012,
		12'h013,
		12'h014,
		12'h015,
		12'h016,
		12'h017,
		12'h018,
		12'h019,
		12'h01a,
		12'h01b,
		12'h01c,
		12'h01d,
		12'h01e,
		12'h01f,
		12'h020,
		12'h021,
		12'h022,
		12'h023,
		12'h024,
		12'h025,
		12'h026,
		12'h027,
		12'h028,
		12'h029,
		12'h02a,
		12'h02b,
		12'h02c,
		12'h02d,
		12'h02e,
		12'h02f,
		12'h030,
		12'h031,
		12'h032,
		12'h033,
		12'h034,
		12'h035,
		12'h036,
		12'h037,
		12'h038,
		12'h039,
		12'h03a,
		12'h03b,
		12'h03c,
		12'h03d,
		12'h03e,
		12'h03f,
		12'h040,
		12'h041,
		12'h042,
		12'h043,
		12'h044,
		12'h045,
		12'h046,
		12'h047,
		12'h048,
		12'h049,
		12'h04a,
		12'h04b,
		12'h04c,
		12'h04d,
		12'h04e,
		12'h04f,
		12'h050,
		12'h051,
		12'h052,
		12'h053,
		12'h054,
		12'h055,
		12'h056,
		12'h057,
		12'h058,
		12'h059,
		12'h05a,
		12'h05b,
		12'h05c,
		12'h05d,
		12'h05e,
		12'h05f,
		12'h060,
		12'h061,
		12'h062,
		12'h063,
		12'h064,
		12'h065,
		12'h066,
		12'h067,
		12'h068,
		12'h069,
		12'h06a,
		12'h06b,
		12'h06c,
		12'h06d,
		12'h06e,
		12'h06f,
		12'h070,
		12'h071,
		12'h072,
		12'h073,
		12'h074,
		12'h075,
		12'h076,
		12'h077,
		12'h078,
		12'h079,
		12'h07a,
		12'h07b,
		12'h07c,
		12'h07d,
		12'h07e,
		12'h07f,
		12'h080,
		12'h081,
		12'h082,
		12'h083,
		12'h084,
		12'h085,
		12'h086,
		12'h087,
		12'h088,
		12'h089,
		12'h08a,
		12'h08b,
		12'h08c,
		12'h08d,
		12'h08e,
		12'h08f,
		12'h090,
		12'h091,
		12'h092,
		12'h093,
		12'h094,
		12'h095,
		12'h096,
		12'h097,
		12'h098,
		12'h099,
		12'h09a,
		12'h09b,
		12'h09c,
		12'h09d,
		12'h09e,
		12'h09f,
		12'h0a0,
		12'h0a1,
		12'h0a2,
		12'h0a3,
		12'h0a4,
		12'h0a5,
		12'h0a6,
		12'h0a7,
		12'h0a8,
		12'h0a9,
		12'h0aa,
		12'h0ab,
		12'h0ac,
		12'h0ad,
		12'h0ae,
		12'h0af,
		12'h0b0,
		12'h0b1,
		12'h0b2,
		12'h0b3,
		12'h0b4,
		12'h0b5,
		12'h0b6,
		12'h0b7,
		12'h0b8,
		12'h0b9,
		12'h0ba,
		12'h0bb,
		12'h0bc,
		12'h0bd,
		12'h0be,
		12'h0bf,
		12'h0c0,
		12'h0c1,
		12'h0c2,
		12'h0c3,
		12'h0c4,
		12'h0c5,
		12'h0c6,
		12'h0c7,
		12'h0c8,
		12'h0c9,
		12'h0ca,
		12'h0cb,
		12'h0cc,
		12'h0cd,
		12'h0ce,
		12'h0cf,
		12'h0d0,
		12'h0d1,
		12'h0d2,
		12'h0d3,
		12'h0d4,
		12'h0d5,
		12'h0d6,
		12'h0d7,
		12'h0d8,
		12'h0d9,
		12'h0da,
		12'h0db,
		12'h0dc,
		12'h0dd,
		12'h0de,
		12'h0df,
		12'h0e0,
		12'h0e1,
		12'h0e2,
		12'h0e3,
		12'h0e4,
		12'h0e5,
		12'h0e6,
		12'h0e7,
		12'h0e8,
		12'h0e9,
		12'h0ea,
		12'h0eb,
		12'h0ec,
		12'h0ed,
		12'h0ee,
		12'h0ef,
		12'h0f0,
		12'h0f1,
		12'h0f2,
		12'h0f3,
		12'h0f4,
		12'h0f5,
		12'h0f6,
		12'h0f7,
		12'h0f8,
		12'h0f9,
		12'h0fa,
		12'h0fb,
		12'h0fc,
		12'h0fd,
		12'h0fe,
		12'h0ff,
		12'h100,
		12'h101,
		12'h102,
		12'h103,
		12'h104,
		12'h105,
		12'h106,
		12'h107,
		12'h108,
		12'h109,
		12'h10a,
		12'h10b,
		12'h10c,
		12'h10d,
		12'h10e,
		12'h10f,
		12'h110,
		12'h111,
		12'h112,
		12'h113,
		12'h114,
		12'h115,
		12'h116,
		12'h117,
		12'h118,
		12'h119,
		12'h11a,
		12'h11b,
		12'h11c,
		12'h11d,
		12'h11e,
		12'h11f,
		12'h120,
		12'h121,
		12'h122,
		12'h123,
		12'h124,
		12'h125,
		12'h126,
		12'h127,
		12'h128,
		12'h129,
		12'h12a,
		12'h12b,
		12'h12c,
		12'h12d,
		12'h12e,
		12'h12f,
		12'h130,
		12'h131,
		12'h132,
		12'h133,
		12'h134,
		12'h135,
		12'h136,
		12'h137,
		12'h138,
		12'h139,
		12'h13a,
		12'h13b,
		12'h13c,
		12'h13d,
		12'h13e,
		12'h13f,
		12'h140,
		12'h141,
		12'h142,
		12'h143,
		12'h144,
		12'h145,
		12'h146,
		12'h147,
		12'h148,
		12'h149,
		12'h14a,
		12'h14b,
		12'h14c,
		12'h14d,
		12'h14e,
		12'h14f,
		12'h150,
		12'h151,
		12'h152,
		12'h153,
		12'h154,
		12'h155,
		12'h156,
		12'h157,
		12'h158,
		12'h159,
		12'h15a,
		12'h15b,
		12'h15c,
		12'h15d,
		12'h15e,
		12'h15f,
		12'h160,
		12'h161,
		12'h162,
		12'h163,
		12'h164,
		12'h165,
		12'h166,
		12'h167,
		12'h168,
		12'h169,
		12'h16a,
		12'h16b,
		12'h16c,
		12'h16d,
		12'h16e,
		12'h16f,
		12'h170,
		12'h171,
		12'h172,
		12'h173,
		12'h174,
		12'h175,
		12'h176,
		12'h177,
		12'h178,
		12'h179,
		12'h17a,
		12'h17b,
		12'h17c,
		12'h17d,
		12'h17e,
		12'h17f,
		12'h180,
		12'h181,
		12'h182,
		12'h183,
		12'h184,
		12'h185,
		12'h186,
		12'h187,
		12'h188,
		12'h189,
		12'h18a,
		12'h18b,
		12'h18c,
		12'h18d,
		12'h18e,
		12'h18f,
		12'h190,
		12'h191,
		12'h192,
		12'h193,
		12'h194,
		12'h195,
		12'h196,
		12'h197,
		12'h198,
		12'h199,
		12'h19a,
		12'h19b,
		12'h19c,
		12'h19d,
		12'h19e,
		12'h19f,
		12'h1a0,
		12'h1a1,
		12'h1a2,
		12'h1a3,
		12'h1a4,
		12'h1a5,
		12'h1a6,
		12'h1a7,
		12'h1a8,
		12'h1a9,
		12'h1aa,
		12'h1ab,
		12'h1ac,
		12'h1ad,
		12'h1ae,
		12'h1af,
		12'h1b0,
		12'h1b1,
		12'h1b2,
		12'h1b3,
		12'h1b4,
		12'h1b5,
		12'h1b6,
		12'h1b7,
		12'h1b8,
		12'h1b9,
		12'h1ba,
		12'h1bb,
		12'h1bc,
		12'h1bd,
		12'h1be,
		12'h1bf,
		12'h1c0,
		12'h1c1,
		12'h1c2,
		12'h1c3,
		12'h1c4,
		12'h1c5,
		12'h1c6,
		12'h1c7,
		12'h1c8,
		12'h1c9,
		12'h1ca,
		12'h1cb,
		12'h1cc,
		12'h1cd,
		12'h1ce,
		12'h1cf,
		12'h1d0,
		12'h1d1,
		12'h1d2,
		12'h1d3,
		12'h1d4,
		12'h1d5,
		12'h1d6,
		12'h1d7,
		12'h1d8,
		12'h1d9,
		12'h1da,
		12'h1db,
		12'h1dc,
		12'h1dd,
		12'h1de,
		12'h1df,
		12'h1e0,
		12'h1e1,
		12'h1e2,
		12'h1e3,
		12'h1e4,
		12'h1e5,
		12'h1e6,
		12'h1e7,
		12'h1e8,
		12'h1e9,
		12'h1ea,
		12'h1eb,
		12'h1ec,
		12'h1ed,
		12'h1ee,
		12'h1ef,
		12'h1f0,
		12'h1f1,
		12'h1f2,
		12'h1f3,
		12'h1f4,
		12'h1f5,
		12'h1f6,
		12'h1f7,
		12'h1f8,
		12'h1f9,
		12'h1fa,
		12'h1fb,
		12'h1fc,
		12'h1fd,
		12'h1fe,
		12'h1ff,
		12'h200,
		12'h201,
		12'h202,
		12'h203,
		12'h204,
		12'h205,
		12'h206,
		12'h207,
		12'h208,
		12'h209,
		12'h20a,
		12'h20b,
		12'h20c,
		12'h20d,
		12'h20e,
		12'h20f,
		12'h210,
		12'h211,
		12'h212,
		12'h213,
		12'h214,
		12'h215,
		12'h216,
		12'h217,
		12'h218,
		12'h219,
		12'h21a,
		12'h21b,
		12'h21c,
		12'h21d,
		12'h21e,
		12'h21f,
		12'h220,
		12'h221,
		12'h222,
		12'h223,
		12'h224,
		12'h225,
		12'h226,
		12'h227,
		12'h228,
		12'h229,
		12'h22a,
		12'h22b,
		12'h22c,
		12'h22d,
		12'h22e,
		12'h22f,
		12'h230,
		12'h231,
		12'h232,
		12'h233,
		12'h234,
		12'h235,
		12'h236,
		12'h237,
		12'h238,
		12'h239,
		12'h23a,
		12'h23b,
		12'h23c,
		12'h23d,
		12'h23e,
		12'h23f,
		12'h240,
		12'h241,
		12'h242,
		12'h243,
		12'h244,
		12'h245,
		12'h246,
		12'h247,
		12'h248,
		12'h249,
		12'h24a,
		12'h24b,
		12'h24c,
		12'h24d,
		12'h24e,
		12'h24f,
		12'h250,
		12'h251,
		12'h252,
		12'h253,
		12'h254,
		12'h255,
		12'h256,
		12'h257,
		12'h258,
		12'h259,
		12'h25a,
		12'h25b,
		12'h25c,
		12'h25d,
		12'h25e,
		12'h25f,
		12'h260,
		12'h261,
		12'h262,
		12'h263,
		12'h264,
		12'h265,
		12'h266,
		12'h267,
		12'h268,
		12'h269,
		12'h26a,
		12'h26b,
		12'h26c,
		12'h26d,
		12'h26e,
		12'h26f,
		12'h270,
		12'h271,
		12'h272,
		12'h273,
		12'h274,
		12'h275,
		12'h276,
		12'h277,
		12'h278,
		12'h279,
		12'h27a,
		12'h27b,
		12'h27c,
		12'h27d,
		12'h27e,
		12'h27f,
		12'h280,
		12'h281,
		12'h282,
		12'h283,
		12'h284,
		12'h285,
		12'h286,
		12'h287,
		12'h288,
		12'h289,
		12'h28a,
		12'h28b,
		12'h28c,
		12'h28d,
		12'h28e,
		12'h28f,
		12'h290,
		12'h291,
		12'h292,
		12'h293,
		12'h294,
		12'h295,
		12'h296,
		12'h297,
		12'h298,
		12'h299,
		12'h29a,
		12'h29b,
		12'h29c,
		12'h29d,
		12'h29e,
		12'h29f,
		12'h2a0,
		12'h2a1,
		12'h2a2,
		12'h2a3,
		12'h2a4,
		12'h2a5,
		12'h2a6,
		12'h2a7,
		12'h2a8,
		12'h2a9,
		12'h2aa,
		12'h2ab,
		12'h2ac,
		12'h2ad,
		12'h2ae,
		12'h2af,
		12'h2b0,
		12'h2b1,
		12'h2b2,
		12'h2b3,
		12'h2b4,
		12'h2b5,
		12'h2b6,
		12'h2b7,
		12'h2b8,
		12'h2b9,
		12'h2ba,
		12'h2bb,
		12'h2bc,
		12'h2bd,
		12'h2be,
		12'h2bf,
		12'h2c0,
		12'h2c1,
		12'h2c2,
		12'h2c3,
		12'h2c4,
		12'h2c5,
		12'h2c6,
		12'h2c7,
		12'h2c8,
		12'h2c9,
		12'h2ca,
		12'h2cb,
		12'h2cc,
		12'h2cd,
		12'h2ce,
		12'h2cf,
		12'h2d0,
		12'h2d1,
		12'h2d2,
		12'h2d3,
		12'h2d4,
		12'h2d5,
		12'h2d6,
		12'h2d7,
		12'h2d8,
		12'h2d9,
		12'h2da,
		12'h2db,
		12'h2dc,
		12'h2dd,
		12'h2de,
		12'h2df,
		12'h2e0,
		12'h2e1,
		12'h2e2,
		12'h2e3,
		12'h2e4,
		12'h2e5,
		12'h2e6,
		12'h2e7,
		12'h2e8,
		12'h2e9,
		12'h2ea,
		12'h2eb,
		12'h2ec,
		12'h2ed,
		12'h2ee,
		12'h2ef,
		12'h2f0,
		12'h2f1,
		12'h2f2,
		12'h2f3,
		12'h2f4,
		12'h2f5,
		12'h2f6,
		12'h2f7,
		12'h2f8,
		12'h2f9,
		12'h2fa,
		12'h2fb,
		12'h2fc,
		12'h2fd,
		12'h2fe,
		12'h2ff,
		12'h300,
		12'h301,
		12'h302,
		12'h303,
		12'h304,
		12'h305,
		12'h306,
		12'h307,
		12'h308,
		12'h309,
		12'h30a,
		12'h30b,
		12'h30c,
		12'h30d,
		12'h30e,
		12'h30f,
		12'h310,
		12'h311,
		12'h312,
		12'h313,
		12'h314,
		12'h315,
		12'h316,
		12'h317,
		12'h318,
		12'h319,
		12'h31a,
		12'h31b,
		12'h31c,
		12'h31d,
		12'h31e,
		12'h31f,
		12'h320,
		12'h321,
		12'h322,
		12'h323,
		12'h324,
		12'h325,
		12'h326,
		12'h327,
		12'h328,
		12'h329,
		12'h32a,
		12'h32b,
		12'h32c,
		12'h32d,
		12'h32e,
		12'h32f,
		12'h330,
		12'h331,
		12'h332,
		12'h333,
		12'h334,
		12'h335,
		12'h336,
		12'h337,
		12'h338,
		12'h339,
		12'h33a,
		12'h33b,
		12'h33c,
		12'h33d,
		12'h33e,
		12'h33f,
		12'h340,
		12'h341,
		12'h342,
		12'h343,
		12'h344,
		12'h345,
		12'h346,
		12'h347,
		12'h348,
		12'h349,
		12'h34a,
		12'h34b,
		12'h34c,
		12'h34d,
		12'h34e,
		12'h34f,
		12'h350,
		12'h351,
		12'h352,
		12'h353,
		12'h354,
		12'h355,
		12'h356,
		12'h357,
		12'h358,
		12'h359,
		12'h35a,
		12'h35b,
		12'h35c,
		12'h35d,
		12'h35e,
		12'h35f,
		12'h360,
		12'h361,
		12'h362,
		12'h363,
		12'h364,
		12'h365,
		12'h366,
		12'h367,
		12'h368,
		12'h369,
		12'h36a,
		12'h36b,
		12'h36c,
		12'h36d,
		12'h36e,
		12'h36f,
		12'h370,
		12'h371,
		12'h372,
		12'h373,
		12'h374,
		12'h375,
		12'h376,
		12'h377,
		12'h378,
		12'h379,
		12'h37a,
		12'h37b,
		12'h37c,
		12'h37d,
		12'h37e,
		12'h37f,
		12'h380,
		12'h381,
		12'h382,
		12'h383,
		12'h384,
		12'h385,
		12'h386,
		12'h387,
		12'h388,
		12'h389,
		12'h38a,
		12'h38b,
		12'h38c,
		12'h38d,
		12'h38e,
		12'h38f,
		12'h390,
		12'h391,
		12'h392,
		12'h393,
		12'h394,
		12'h395,
		12'h396,
		12'h397,
		12'h398,
		12'h399,
		12'h39a,
		12'h39b,
		12'h39c,
		12'h39d,
		12'h39e,
		12'h39f,
		12'h3a0,
		12'h3a1,
		12'h3a2,
		12'h3a3,
		12'h3a4,
		12'h3a5,
		12'h3a6,
		12'h3a7,
		12'h3a8,
		12'h3a9,
		12'h3aa,
		12'h3ab,
		12'h3ac,
		12'h3ad,
		12'h3ae,
		12'h3af,
		12'h3b0,
		12'h3b1,
		12'h3b2,
		12'h3b3,
		12'h3b4,
		12'h3b5,
		12'h3b6,
		12'h3b7,
		12'h3b8,
		12'h3b9,
		12'h3ba,
		12'h3bb,
		12'h3bc,
		12'h3bd,
		12'h3be,
		12'h3bf,
		12'h3c0,
		12'h3c1,
		12'h3c2,
		12'h3c3,
		12'h3c4,
		12'h3c5,
		12'h3c6,
		12'h3c7,
		12'h3c8,
		12'h3c9,
		12'h3ca,
		12'h3cb,
		12'h3cc,
		12'h3cd,
		12'h3ce,
		12'h3cf,
		12'h3d0,
		12'h3d1,
		12'h3d2,
		12'h3d3,
		12'h3d4,
		12'h3d5,
		12'h3d6,
		12'h3d7,
		12'h3d8,
		12'h3d9,
		12'h3da,
		12'h3db,
		12'h3dc,
		12'h3dd,
		12'h3de,
		12'h3df,
		12'h3e0,
		12'h3e1,
		12'h3e2,
		12'h3e3,
		12'h3e4,
		12'h3e5,
		12'h3e6,
		12'h3e7,
		12'h3e8,
		12'h3e9,
		12'h3ea,
		12'h3eb,
		12'h3ec,
		12'h3ed,
		12'h3ee,
		12'h3ef,
		12'h3f0,
		12'h3f1,
		12'h3f2,
		12'h3f3,
		12'h3f4,
		12'h3f5,
		12'h3f6,
		12'h3f7,
		12'h3f8,
		12'h3f9,
		12'h3fa,
		12'h3fb,
		12'h3fc,
		12'h3fd,
		12'h3fe,
		12'h3ff,
		12'h400,
		12'h401,
		12'h402,
		12'h403,
		12'h404,
		12'h405,
		12'h406,
		12'h407,
		12'h408,
		12'h409,
		12'h40a,
		12'h40b,
		12'h40c,
		12'h40d,
		12'h40e,
		12'h40f,
		12'h410,
		12'h411,
		12'h412,
		12'h413,
		12'h414,
		12'h415,
		12'h416,
		12'h417,
		12'h418,
		12'h419,
		12'h41a,
		12'h41b,
		12'h41c,
		12'h41d,
		12'h41e,
		12'h41f,
		12'h420,
		12'h421,
		12'h422,
		12'h423,
		12'h424,
		12'h425,
		12'h426,
		12'h427,
		12'h428,
		12'h429,
		12'h42a,
		12'h42b,
		12'h42c,
		12'h42d,
		12'h42e,
		12'h42f,
		12'h430,
		12'h431,
		12'h432,
		12'h433,
		12'h434,
		12'h435,
		12'h436,
		12'h437,
		12'h438,
		12'h439,
		12'h43a,
		12'h43b,
		12'h43c,
		12'h43d,
		12'h43e,
		12'h43f,
		12'h440,
		12'h441,
		12'h442,
		12'h443,
		12'h444,
		12'h445,
		12'h446,
		12'h447,
		12'h448,
		12'h449,
		12'h44a,
		12'h44b,
		12'h44c,
		12'h44d,
		12'h44e,
		12'h44f,
		12'h450,
		12'h451,
		12'h452,
		12'h453,
		12'h454,
		12'h455,
		12'h456,
		12'h457,
		12'h458,
		12'h459,
		12'h45a,
		12'h45b,
		12'h45c,
		12'h45d,
		12'h45e,
		12'h45f,
		12'h460,
		12'h461,
		12'h462,
		12'h463,
		12'h464,
		12'h465,
		12'h466,
		12'h467,
		12'h468,
		12'h469,
		12'h46a,
		12'h46b,
		12'h46c,
		12'h46d,
		12'h46e,
		12'h46f,
		12'h470,
		12'h471,
		12'h472,
		12'h473,
		12'h474,
		12'h475,
		12'h476,
		12'h477,
		12'h478,
		12'h479,
		12'h47a,
		12'h47b,
		12'h47c,
		12'h47d,
		12'h47e,
		12'h47f,
		12'h480,
		12'h481,
		12'h482,
		12'h483,
		12'h484,
		12'h485,
		12'h486,
		12'h487,
		12'h488,
		12'h489,
		12'h48a,
		12'h48b,
		12'h48c,
		12'h48d,
		12'h48e,
		12'h48f,
		12'h490,
		12'h491,
		12'h492,
		12'h493,
		12'h494,
		12'h495,
		12'h496,
		12'h497,
		12'h498,
		12'h499,
		12'h49a,
		12'h49b,
		12'h49c,
		12'h49d,
		12'h49e,
		12'h49f,
		12'h4a0,
		12'h4a1,
		12'h4a2,
		12'h4a3,
		12'h4a4,
		12'h4a5,
		12'h4a6,
		12'h4a7,
		12'h4a8,
		12'h4a9,
		12'h4aa,
		12'h4ab,
		12'h4ac,
		12'h4ad,
		12'h4ae,
		12'h4af,
		12'h4b0,
		12'h4b1,
		12'h4b2,
		12'h4b3,
		12'h4b4,
		12'h4b5,
		12'h4b6,
		12'h4b7,
		12'h4b8,
		12'h4b9,
		12'h4ba,
		12'h4bb,
		12'h4bc,
		12'h4bd,
		12'h4be,
		12'h4bf,
		12'h4c0,
		12'h4c1,
		12'h4c2,
		12'h4c3,
		12'h4c4,
		12'h4c5,
		12'h4c6,
		12'h4c7,
		12'h4c8,
		12'h4c9,
		12'h4ca,
		12'h4cb,
		12'h4cc,
		12'h4cd,
		12'h4ce,
		12'h4cf,
		12'h4d0,
		12'h4d1,
		12'h4d2,
		12'h4d3,
		12'h4d4,
		12'h4d5,
		12'h4d6,
		12'h4d7,
		12'h4d8,
		12'h4d9,
		12'h4da,
		12'h4db,
		12'h4dc,
		12'h4dd,
		12'h4de,
		12'h4df,
		12'h4e0,
		12'h4e1,
		12'h4e2,
		12'h4e3,
		12'h4e4,
		12'h4e5,
		12'h4e6,
		12'h4e7,
		12'h4e8,
		12'h4e9,
		12'h4ea,
		12'h4eb,
		12'h4ec,
		12'h4ed,
		12'h4ee,
		12'h4ef,
		12'h4f0,
		12'h4f1,
		12'h4f2,
		12'h4f3,
		12'h4f4,
		12'h4f5,
		12'h4f6,
		12'h4f7,
		12'h4f8,
		12'h4f9,
		12'h4fa,
		12'h4fb,
		12'h4fc,
		12'h4fd,
		12'h4fe,
		12'h4ff,
		12'h500,
		12'h501,
		12'h502,
		12'h503,
		12'h504,
		12'h505,
		12'h506,
		12'h507,
		12'h508,
		12'h509,
		12'h50a,
		12'h50b,
		12'h50c,
		12'h50d,
		12'h50e,
		12'h50f,
		12'h510,
		12'h511,
		12'h512,
		12'h513,
		12'h514,
		12'h515,
		12'h516,
		12'h517,
		12'h518,
		12'h519,
		12'h51a,
		12'h51b,
		12'h51c,
		12'h51d,
		12'h51e,
		12'h51f,
		12'h520,
		12'h521,
		12'h522,
		12'h523,
		12'h524,
		12'h525,
		12'h526,
		12'h527,
		12'h528,
		12'h529,
		12'h52a,
		12'h52b,
		12'h52c,
		12'h52d,
		12'h52e,
		12'h52f,
		12'h530,
		12'h531,
		12'h532,
		12'h533,
		12'h534,
		12'h535,
		12'h536,
		12'h537,
		12'h538,
		12'h539,
		12'h53a,
		12'h53b,
		12'h53c,
		12'h53d,
		12'h53e,
		12'h53f,
		12'h540,
		12'h541,
		12'h542,
		12'h543,
		12'h544,
		12'h545,
		12'h546,
		12'h547,
		12'h548,
		12'h549,
		12'h54a,
		12'h54b,
		12'h54c,
		12'h54d,
		12'h54e,
		12'h54f,
		12'h550,
		12'h551,
		12'h552,
		12'h553,
		12'h554,
		12'h555,
		12'h556,
		12'h557,
		12'h558,
		12'h559,
		12'h55a,
		12'h55b,
		12'h55c,
		12'h55d,
		12'h55e,
		12'h55f,
		12'h560,
		12'h561,
		12'h562,
		12'h563,
		12'h564,
		12'h565,
		12'h566,
		12'h567,
		12'h568,
		12'h569,
		12'h56a,
		12'h56b,
		12'h56c,
		12'h56d,
		12'h56e,
		12'h56f,
		12'h570,
		12'h571,
		12'h572,
		12'h573,
		12'h574,
		12'h575,
		12'h576,
		12'h577,
		12'h578,
		12'h579,
		12'h57a,
		12'h57b,
		12'h57c,
		12'h57d,
		12'h57e,
		12'h57f,
		12'h580,
		12'h581,
		12'h582,
		12'h583,
		12'h584,
		12'h585,
		12'h586,
		12'h587,
		12'h588,
		12'h589,
		12'h58a,
		12'h58b,
		12'h58c,
		12'h58d,
		12'h58e,
		12'h58f,
		12'h590,
		12'h591,
		12'h592,
		12'h593,
		12'h594,
		12'h595,
		12'h596,
		12'h597,
		12'h598,
		12'h599,
		12'h59a,
		12'h59b,
		12'h59c,
		12'h59d,
		12'h59e,
		12'h59f,
		12'h5a0,
		12'h5a1,
		12'h5a2,
		12'h5a3,
		12'h5a4,
		12'h5a5,
		12'h5a6,
		12'h5a7,
		12'h5a8,
		12'h5a9,
		12'h5aa,
		12'h5ab,
		12'h5ac,
		12'h5ad,
		12'h5ae,
		12'h5af,
		12'h5b0,
		12'h5b1,
		12'h5b2,
		12'h5b3,
		12'h5b4,
		12'h5b5,
		12'h5b6,
		12'h5b7,
		12'h5b8,
		12'h5b9,
		12'h5ba,
		12'h5bb,
		12'h5bc,
		12'h5bd,
		12'h5be,
		12'h5bf,
		12'h5c0,
		12'h5c1,
		12'h5c2,
		12'h5c3,
		12'h5c4,
		12'h5c5,
		12'h5c6,
		12'h5c7,
		12'h5c8,
		12'h5c9,
		12'h5ca,
		12'h5cb,
		12'h5cc,
		12'h5cd,
		12'h5ce,
		12'h5cf,
		12'h5d0,
		12'h5d1,
		12'h5d2,
		12'h5d3,
		12'h5d4,
		12'h5d5,
		12'h5d6,
		12'h5d7,
		12'h5d8,
		12'h5d9,
		12'h5da,
		12'h5db,
		12'h5dc,
		12'h5dd,
		12'h5de,
		12'h5df,
		12'h5e0,
		12'h5e1,
		12'h5e2,
		12'h5e3,
		12'h5e4,
		12'h5e5,
		12'h5e6,
		12'h5e7,
		12'h5e8,
		12'h5e9,
		12'h5ea,
		12'h5eb,
		12'h5ec,
		12'h5ed,
		12'h5ee,
		12'h5ef,
		12'h5f0,
		12'h5f1,
		12'h5f2,
		12'h5f3,
		12'h5f4,
		12'h5f5,
		12'h5f6,
		12'h5f7,
		12'h5f8,
		12'h5f9,
		12'h5fa,
		12'h5fb,
		12'h5fc,
		12'h5fd,
		12'h5fe,
		12'h5ff,
		12'h600,
		12'h601,
		12'h602,
		12'h603,
		12'h604,
		12'h605,
		12'h606,
		12'h607,
		12'h608,
		12'h609,
		12'h60a,
		12'h60b,
		12'h60c,
		12'h60d,
		12'h60e,
		12'h60f,
		12'h610,
		12'h611,
		12'h612,
		12'h613,
		12'h614,
		12'h615,
		12'h616,
		12'h617,
		12'h618,
		12'h619,
		12'h61a,
		12'h61b,
		12'h61c,
		12'h61d,
		12'h61e,
		12'h61f,
		12'h620,
		12'h621,
		12'h622,
		12'h623,
		12'h624,
		12'h625,
		12'h626,
		12'h627,
		12'h628,
		12'h629,
		12'h62a,
		12'h62b,
		12'h62c,
		12'h62d,
		12'h62e,
		12'h62f,
		12'h630,
		12'h631,
		12'h632,
		12'h633,
		12'h634,
		12'h635,
		12'h636,
		12'h637,
		12'h638,
		12'h639,
		12'h63a,
		12'h63b,
		12'h63c,
		12'h63d,
		12'h63e,
		12'h63f,
		12'h640,
		12'h641,
		12'h642,
		12'h643,
		12'h644,
		12'h645,
		12'h646,
		12'h647,
		12'h648,
		12'h649,
		12'h64a,
		12'h64b,
		12'h64c,
		12'h64d,
		12'h64e,
		12'h64f,
		12'h650,
		12'h651,
		12'h652,
		12'h653,
		12'h654,
		12'h655,
		12'h656,
		12'h657,
		12'h658,
		12'h659,
		12'h65a,
		12'h65b,
		12'h65c,
		12'h65d,
		12'h65e,
		12'h65f,
		12'h660,
		12'h661,
		12'h662,
		12'h663,
		12'h664,
		12'h665,
		12'h666,
		12'h667,
		12'h668,
		12'h669,
		12'h66a,
		12'h66b,
		12'h66c,
		12'h66d,
		12'h66e,
		12'h66f,
		12'h670,
		12'h671,
		12'h672,
		12'h673,
		12'h674,
		12'h675,
		12'h676,
		12'h677,
		12'h678,
		12'h679,
		12'h67a,
		12'h67b,
		12'h67c,
		12'h67d,
		12'h67e,
		12'h67f,
		12'h680,
		12'h681,
		12'h682,
		12'h683,
		12'h684,
		12'h685,
		12'h686,
		12'h687,
		12'h688,
		12'h689,
		12'h68a,
		12'h68b,
		12'h68c,
		12'h68d,
		12'h68e,
		12'h68f,
		12'h690,
		12'h691,
		12'h692,
		12'h693,
		12'h694,
		12'h695,
		12'h696,
		12'h697,
		12'h698,
		12'h699,
		12'h69a,
		12'h69b,
		12'h69c,
		12'h69d,
		12'h69e,
		12'h69f,
		12'h6a0,
		12'h6a1,
		12'h6a2,
		12'h6a3,
		12'h6a4,
		12'h6a5,
		12'h6a6,
		12'h6a7,
		12'h6a8,
		12'h6a9,
		12'h6aa,
		12'h6ab,
		12'h6ac,
		12'h6ad,
		12'h6ae,
		12'h6af,
		12'h6b0,
		12'h6b1,
		12'h6b2,
		12'h6b3,
		12'h6b4,
		12'h6b5,
		12'h6b6,
		12'h6b7,
		12'h6b8,
		12'h6b9,
		12'h6ba,
		12'h6bb,
		12'h6bc,
		12'h6bd,
		12'h6be,
		12'h6bf,
		12'h6c0,
		12'h6c1,
		12'h6c2,
		12'h6c3,
		12'h6c4,
		12'h6c5,
		12'h6c6,
		12'h6c7,
		12'h6c8,
		12'h6c9,
		12'h6ca,
		12'h6cb,
		12'h6cc,
		12'h6cd,
		12'h6ce,
		12'h6cf,
		12'h6d0,
		12'h6d1,
		12'h6d2,
		12'h6d3,
		12'h6d4,
		12'h6d5,
		12'h6d6,
		12'h6d7,
		12'h6d8,
		12'h6d9,
		12'h6da,
		12'h6db,
		12'h6dc,
		12'h6dd,
		12'h6de,
		12'h6df,
		12'h6e0,
		12'h6e1,
		12'h6e2,
		12'h6e3,
		12'h6e4,
		12'h6e5,
		12'h6e6,
		12'h6e7,
		12'h6e8,
		12'h6e9,
		12'h6ea,
		12'h6eb,
		12'h6ec,
		12'h6ed,
		12'h6ee,
		12'h6ef,
		12'h6f0,
		12'h6f1,
		12'h6f2,
		12'h6f3,
		12'h6f4,
		12'h6f5,
		12'h6f6,
		12'h6f7,
		12'h6f8,
		12'h6f9,
		12'h6fa,
		12'h6fb,
		12'h6fc,
		12'h6fd,
		12'h6fe,
		12'h6ff,
		12'h700,
		12'h701,
		12'h702,
		12'h703,
		12'h704,
		12'h705,
		12'h706,
		12'h707,
		12'h708,
		12'h709,
		12'h70a,
		12'h70b,
		12'h70c,
		12'h70d,
		12'h70e,
		12'h70f,
		12'h710,
		12'h711,
		12'h712,
		12'h713,
		12'h714,
		12'h715,
		12'h716,
		12'h717,
		12'h718,
		12'h719,
		12'h71a,
		12'h71b,
		12'h71c,
		12'h71d,
		12'h71e,
		12'h71f,
		12'h720,
		12'h721,
		12'h722,
		12'h723,
		12'h724,
		12'h725,
		12'h726,
		12'h727,
		12'h728,
		12'h729,
		12'h72a,
		12'h72b,
		12'h72c,
		12'h72d,
		12'h72e,
		12'h72f,
		12'h730,
		12'h731,
		12'h732,
		12'h733,
		12'h734,
		12'h735,
		12'h736,
		12'h737,
		12'h738,
		12'h739,
		12'h73a,
		12'h73b,
		12'h73c,
		12'h73d,
		12'h73e,
		12'h73f,
		12'h740,
		12'h741,
		12'h742,
		12'h743,
		12'h744,
		12'h745,
		12'h746,
		12'h747,
		12'h748,
		12'h749,
		12'h74a,
		12'h74b,
		12'h74c,
		12'h74d,
		12'h74e,
		12'h74f,
		12'h750,
		12'h751,
		12'h752,
		12'h753,
		12'h754,
		12'h755,
		12'h756,
		12'h757,
		12'h758,
		12'h759,
		12'h75a,
		12'h75b,
		12'h75c,
		12'h75d,
		12'h75e,
		12'h75f,
		12'h760,
		12'h761,
		12'h762,
		12'h763,
		12'h764,
		12'h765,
		12'h766,
		12'h767,
		12'h768,
		12'h769,
		12'h76a,
		12'h76b,
		12'h76c,
		12'h76d,
		12'h76e,
		12'h76f,
		12'h770,
		12'h771,
		12'h772,
		12'h773,
		12'h774,
		12'h775,
		12'h776,
		12'h777,
		12'h778,
		12'h779,
		12'h77a,
		12'h77b,
		12'h77c,
		12'h77d,
		12'h77e,
		12'h77f,
		12'h780,
		12'h781,
		12'h782,
		12'h783,
		12'h784,
		12'h785,
		12'h786,
		12'h787,
		12'h788,
		12'h789,
		12'h78a,
		12'h78b,
		12'h78c,
		12'h78d,
		12'h78e,
		12'h78f,
		12'h790,
		12'h791,
		12'h792,
		12'h793,
		12'h794,
		12'h795,
		12'h796,
		12'h797,
		12'h798,
		12'h799,
		12'h79a,
		12'h79b,
		12'h79c,
		12'h79d,
		12'h79e,
		12'h79f,
		12'h7a0,
		12'h7a1,
		12'h7a2,
		12'h7a3,
		12'h7a4,
		12'h7a5,
		12'h7a6,
		12'h7a7,
		12'h7a8,
		12'h7a9,
		12'h7aa,
		12'h7ab,
		12'h7ac,
		12'h7ad,
		12'h7ae,
		12'h7af,
		12'h7b0,
		12'h7b1,
		12'h7b2,
		12'h7b3,
		12'h7b4,
		12'h7b5,
		12'h7b6,
		12'h7b7,
		12'h7b8,
		12'h7b9,
		12'h7ba,
		12'h7bb,
		12'h7bc,
		12'h7bd,
		12'h7be,
		12'h7bf,
		12'h7c0,
		12'h7c1,
		12'h7c2,
		12'h7c3,
		12'h7c4,
		12'h7c5,
		12'h7c6,
		12'h7c7,
		12'h7c8,
		12'h7c9,
		12'h7ca,
		12'h7cb,
		12'h7cc,
		12'h7cd,
		12'h7ce,
		12'h7cf,
		12'h7d0,
		12'h7d1,
		12'h7d2,
		12'h7d3,
		12'h7d4,
		12'h7d5,
		12'h7d6,
		12'h7d7,
		12'h7d8,
		12'h7d9,
		12'h7da,
		12'h7db,
		12'h7dc,
		12'h7dd,
		12'h7de,
		12'h7df,
		12'h7e0,
		12'h7e1,
		12'h7e2,
		12'h7e3,
		12'h7e4,
		12'h7e5,
		12'h7e6,
		12'h7e7,
		12'h7e8,
		12'h7e9,
		12'h7ea,
		12'h7eb,
		12'h7ec,
		12'h7ed,
		12'h7ee,
		12'h7ef,
		12'h7f0,
		12'h7f1,
		12'h7f2,
		12'h7f3,
		12'h7f4,
		12'h7f5,
		12'h7f6,
		12'h7f7,
		12'h7f8,
		12'h7f9,
		12'h7fa,
		12'h7fb,
		12'h7fc,
		12'h7fd,
		12'h7fe,
		12'h7ff,
		12'h800,
		12'h801,
		12'h802,
		12'h803,
		12'h804,
		12'h805,
		12'h806,
		12'h807,
		12'h808,
		12'h809,
		12'h80a,
		12'h80b,
		12'h80c,
		12'h80d,
		12'h80e,
		12'h80f,
		12'h810,
		12'h811,
		12'h812,
		12'h813,
		12'h814,
		12'h815,
		12'h816,
		12'h817,
		12'h818,
		12'h819,
		12'h81a,
		12'h81b,
		12'h81c,
		12'h81d,
		12'h81e,
		12'h81f,
		12'h820,
		12'h821,
		12'h822,
		12'h823,
		12'h824,
		12'h825,
		12'h826,
		12'h827,
		12'h828,
		12'h829,
		12'h82a,
		12'h82b,
		12'h82c,
		12'h82d,
		12'h82e,
		12'h82f,
		12'h830,
		12'h831,
		12'h832,
		12'h833,
		12'h834,
		12'h835,
		12'h836,
		12'h837,
		12'h838,
		12'h839,
		12'h83a,
		12'h83b,
		12'h83c,
		12'h83d,
		12'h83e,
		12'h83f,
		12'h840,
		12'h841,
		12'h842,
		12'h843,
		12'h844,
		12'h845,
		12'h846,
		12'h847,
		12'h848,
		12'h849,
		12'h84a,
		12'h84b,
		12'h84c,
		12'h84d,
		12'h84e,
		12'h84f,
		12'h850,
		12'h851,
		12'h852,
		12'h853,
		12'h854,
		12'h855,
		12'h856,
		12'h857,
		12'h858,
		12'h859,
		12'h85a,
		12'h85b,
		12'h85c,
		12'h85d,
		12'h85e,
		12'h85f,
		12'h860,
		12'h861,
		12'h862,
		12'h863,
		12'h864,
		12'h865,
		12'h866,
		12'h867,
		12'h868,
		12'h869,
		12'h86a,
		12'h86b,
		12'h86c,
		12'h86d,
		12'h86e,
		12'h86f,
		12'h870,
		12'h871,
		12'h872,
		12'h873,
		12'h874,
		12'h875,
		12'h876,
		12'h877,
		12'h878,
		12'h879,
		12'h87a,
		12'h87b,
		12'h87c,
		12'h87d,
		12'h87e,
		12'h87f,
		12'h880,
		12'h881,
		12'h882,
		12'h883,
		12'h884,
		12'h885,
		12'h886,
		12'h887,
		12'h888,
		12'h889,
		12'h88a,
		12'h88b,
		12'h88c,
		12'h88d,
		12'h88e,
		12'h88f,
		12'h890,
		12'h891,
		12'h892,
		12'h893,
		12'h894,
		12'h895,
		12'h896,
		12'h897,
		12'h898,
		12'h899,
		12'h89a,
		12'h89b,
		12'h89c,
		12'h89d,
		12'h89e,
		12'h89f,
		12'h8a0,
		12'h8a1,
		12'h8a2,
		12'h8a3,
		12'h8a4,
		12'h8a5,
		12'h8a6,
		12'h8a7,
		12'h8a8,
		12'h8a9,
		12'h8aa,
		12'h8ab,
		12'h8ac,
		12'h8ad,
		12'h8ae,
		12'h8af,
		12'h8b0,
		12'h8b1,
		12'h8b2,
		12'h8b3,
		12'h8b4,
		12'h8b5,
		12'h8b6,
		12'h8b7,
		12'h8b8,
		12'h8b9,
		12'h8ba,
		12'h8bb,
		12'h8bc,
		12'h8bd,
		12'h8be,
		12'h8bf,
		12'h8c0,
		12'h8c1,
		12'h8c2,
		12'h8c3,
		12'h8c4,
		12'h8c5,
		12'h8c6,
		12'h8c7,
		12'h8c8,
		12'h8c9,
		12'h8ca,
		12'h8cb,
		12'h8cc,
		12'h8cd,
		12'h8ce,
		12'h8cf,
		12'h8d0,
		12'h8d1,
		12'h8d2,
		12'h8d3,
		12'h8d4,
		12'h8d5,
		12'h8d6,
		12'h8d7,
		12'h8d8,
		12'h8d9,
		12'h8da,
		12'h8db,
		12'h8dc,
		12'h8dd,
		12'h8de,
		12'h8df,
		12'h8e0,
		12'h8e1,
		12'h8e2,
		12'h8e3,
		12'h8e4,
		12'h8e5,
		12'h8e6,
		12'h8e7,
		12'h8e8,
		12'h8e9,
		12'h8ea,
		12'h8eb,
		12'h8ec,
		12'h8ed,
		12'h8ee,
		12'h8ef,
		12'h8f0,
		12'h8f1,
		12'h8f2,
		12'h8f3,
		12'h8f4,
		12'h8f5,
		12'h8f6,
		12'h8f7,
		12'h8f8,
		12'h8f9,
		12'h8fa,
		12'h8fb,
		12'h8fc,
		12'h8fd,
		12'h8fe,
		12'h8ff,
		12'h900,
		12'h901,
		12'h902,
		12'h903,
		12'h904,
		12'h905,
		12'h906,
		12'h907,
		12'h908,
		12'h909,
		12'h90a,
		12'h90b,
		12'h90c,
		12'h90d,
		12'h90e,
		12'h90f,
		12'h910,
		12'h911,
		12'h912,
		12'h913,
		12'h914,
		12'h915,
		12'h916,
		12'h917,
		12'h918,
		12'h919,
		12'h91a,
		12'h91b,
		12'h91c,
		12'h91d,
		12'h91e,
		12'h91f,
		12'h920,
		12'h921,
		12'h922,
		12'h923,
		12'h924,
		12'h925,
		12'h926,
		12'h927,
		12'h928,
		12'h929,
		12'h92a,
		12'h92b,
		12'h92c,
		12'h92d,
		12'h92e,
		12'h92f,
		12'h930,
		12'h931,
		12'h932,
		12'h933,
		12'h934,
		12'h935,
		12'h936,
		12'h937,
		12'h938,
		12'h939,
		12'h93a,
		12'h93b,
		12'h93c,
		12'h93d,
		12'h93e,
		12'h93f,
		12'h940,
		12'h941,
		12'h942,
		12'h943,
		12'h944,
		12'h945,
		12'h946,
		12'h947,
		12'h948,
		12'h949,
		12'h94a,
		12'h94b,
		12'h94c,
		12'h94d,
		12'h94e,
		12'h94f,
		12'h950,
		12'h951,
		12'h952,
		12'h953,
		12'h954,
		12'h955,
		12'h956,
		12'h957,
		12'h958,
		12'h959,
		12'h95a,
		12'h95b,
		12'h95c,
		12'h95d,
		12'h95e,
		12'h95f,
		12'h960,
		12'h961,
		12'h962,
		12'h963,
		12'h964,
		12'h965,
		12'h966,
		12'h967,
		12'h968,
		12'h969,
		12'h96a,
		12'h96b,
		12'h96c,
		12'h96d,
		12'h96e,
		12'h96f,
		12'h970,
		12'h971,
		12'h972,
		12'h973,
		12'h974,
		12'h975,
		12'h976,
		12'h977,
		12'h978,
		12'h979,
		12'h97a,
		12'h97b,
		12'h97c,
		12'h97d,
		12'h97e,
		12'h97f,
		12'h980,
		12'h981,
		12'h982,
		12'h983,
		12'h984,
		12'h985,
		12'h986,
		12'h987,
		12'h988,
		12'h989,
		12'h98a,
		12'h98b,
		12'h98c,
		12'h98d,
		12'h98e,
		12'h98f,
		12'h990,
		12'h991,
		12'h992,
		12'h993,
		12'h994,
		12'h995,
		12'h996,
		12'h997,
		12'h998,
		12'h999,
		12'h99a,
		12'h99b,
		12'h99c,
		12'h99d,
		12'h99e,
		12'h99f,
		12'h9a0,
		12'h9a1,
		12'h9a2,
		12'h9a3,
		12'h9a4,
		12'h9a5,
		12'h9a6,
		12'h9a7,
		12'h9a8,
		12'h9a9,
		12'h9aa,
		12'h9ab,
		12'h9ac,
		12'h9ad,
		12'h9ae,
		12'h9af,
		12'h9b0,
		12'h9b1,
		12'h9b2,
		12'h9b3,
		12'h9b4,
		12'h9b5,
		12'h9b6,
		12'h9b7,
		12'h9b8,
		12'h9b9,
		12'h9ba,
		12'h9bb,
		12'h9bc,
		12'h9bd,
		12'h9be,
		12'h9bf,
		12'h9c0,
		12'h9c1,
		12'h9c2,
		12'h9c3

	
	};

	assign addr = ROM[ycoord][xcoord];
endmodule